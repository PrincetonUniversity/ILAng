module GB(
arg_0_TREADY,
arg_1_TDATA,
arg_1_TVALID,
RAM_w,
RAM_x,
RAM_y,
arg_0_TDATA,
arg_0_TVALID,
arg_1_TREADY,
cur_pix,
pre_pix,
proc_in,
st_ready,
stencil_0,
stencil_1,
stencil_2,
stencil_3,
stencil_4,
stencil_5,
stencil_6,
stencil_7,
stencil_8,
clk,rst,
step
);
input            arg_0_TREADY;
input      [7:0] arg_1_TDATA;
input            arg_1_TVALID;
input clk;
input rst;
input step;
output      [2:0] RAM_w;
output      [8:0] RAM_x;
output      [9:0] RAM_y;
output      [7:0] arg_0_TDATA;
output            arg_0_TVALID;
output            arg_1_TREADY;
output      [7:0] cur_pix;
output      [7:0] pre_pix;
output    [647:0] proc_in;
output            st_ready;
output     [71:0] stencil_0;
output     [71:0] stencil_1;
output     [71:0] stencil_2;
output     [71:0] stencil_3;
output     [71:0] stencil_4;
output     [71:0] stencil_5;
output     [71:0] stencil_6;
output     [71:0] stencil_7;
output     [71:0] stencil_8;
reg      [2:0] RAM_w;
reg      [8:0] RAM_x;
reg      [9:0] RAM_y;
reg      [7:0] arg_0_TDATA;
reg            arg_0_TVALID;
reg            arg_1_TREADY;
reg      [7:0] cur_pix;
reg      [7:0] pre_pix;
reg    [647:0] proc_in;
reg            st_ready;
reg     [71:0] stencil_0;
reg     [71:0] stencil_1;
reg     [71:0] stencil_2;
reg     [71:0] stencil_3;
reg     [71:0] stencil_4;
reg     [71:0] stencil_5;
reg     [71:0] stencil_6;
reg     [71:0] stencil_7;
reg     [71:0] stencil_8;
wire            arg_0_TREADY;
wire      [7:0] arg_1_TDATA;
wire            arg_1_TVALID;
wire            n0;
wire            n1;
wire            n2;
wire            n3;
wire            n4;
wire            n5;
wire            n6;
wire            n7;
wire            n8;
wire            n9;
wire            n10;
wire            n11;
wire            n12;
wire            n13;
wire            n14;
wire            n15;
wire            n16;
wire            n17;
wire            n18;
wire      [2:0] n19;
wire      [2:0] n20;
wire      [2:0] n21;
wire            n22;
wire            n23;
wire            n24;
wire            n25;
wire            n26;
wire      [2:0] n27;
wire      [2:0] n28;
wire      [2:0] n29;
wire      [2:0] n30;
wire      [8:0] n31;
wire      [8:0] n32;
wire      [8:0] n33;
wire      [8:0] n34;
wire      [8:0] n35;
wire      [8:0] n36;
wire            n37;
wire      [9:0] n38;
wire      [9:0] n39;
wire      [9:0] n40;
wire      [9:0] n41;
wire      [9:0] n42;
wire      [9:0] n43;
wire      [9:0] n44;
wire            n45;
wire            n46;
wire            n47;
wire      [7:0] n48;
wire      [7:0] n49;
wire      [7:0] n50;
wire      [7:0] n51;
wire      [7:0] n52;
wire      [7:0] n53;
wire      [7:0] n54;
wire      [7:0] n55;
wire      [7:0] n56;
wire     [15:0] n57;
wire     [23:0] n58;
wire     [31:0] n59;
wire     [39:0] n60;
wire     [47:0] n61;
wire     [55:0] n62;
wire     [63:0] n63;
wire     [71:0] n64;
wire      [7:0] n65;
wire      [7:0] n66;
wire      [7:0] n67;
wire      [7:0] n68;
wire      [7:0] n69;
wire      [7:0] n70;
wire      [7:0] n71;
wire      [7:0] n72;
wire      [7:0] n73;
wire     [15:0] n74;
wire     [23:0] n75;
wire     [31:0] n76;
wire     [39:0] n77;
wire     [47:0] n78;
wire     [55:0] n79;
wire     [63:0] n80;
wire     [71:0] n81;
wire      [7:0] n82;
wire      [7:0] n83;
wire      [7:0] n84;
wire      [7:0] n85;
wire      [7:0] n86;
wire      [7:0] n87;
wire      [7:0] n88;
wire      [7:0] n89;
wire      [7:0] n90;
wire     [15:0] n91;
wire     [23:0] n92;
wire     [31:0] n93;
wire     [39:0] n94;
wire     [47:0] n95;
wire     [55:0] n96;
wire     [63:0] n97;
wire     [71:0] n98;
wire      [7:0] n99;
wire      [7:0] n100;
wire      [7:0] n101;
wire      [7:0] n102;
wire      [7:0] n103;
wire      [7:0] n104;
wire      [7:0] n105;
wire      [7:0] n106;
wire      [7:0] n107;
wire     [15:0] n108;
wire     [23:0] n109;
wire     [31:0] n110;
wire     [39:0] n111;
wire     [47:0] n112;
wire     [55:0] n113;
wire     [63:0] n114;
wire     [71:0] n115;
wire      [7:0] n116;
wire      [7:0] n117;
wire      [7:0] n118;
wire      [7:0] n119;
wire      [7:0] n120;
wire      [7:0] n121;
wire      [7:0] n122;
wire      [7:0] n123;
wire      [7:0] n124;
wire     [15:0] n125;
wire     [23:0] n126;
wire     [31:0] n127;
wire     [39:0] n128;
wire     [47:0] n129;
wire     [55:0] n130;
wire     [63:0] n131;
wire     [71:0] n132;
wire      [7:0] n133;
wire      [7:0] n134;
wire      [7:0] n135;
wire      [7:0] n136;
wire      [7:0] n137;
wire      [7:0] n138;
wire      [7:0] n139;
wire      [7:0] n140;
wire      [7:0] n141;
wire     [15:0] n142;
wire     [23:0] n143;
wire     [31:0] n144;
wire     [39:0] n145;
wire     [47:0] n146;
wire     [55:0] n147;
wire     [63:0] n148;
wire     [71:0] n149;
wire      [7:0] n150;
wire      [7:0] n151;
wire      [7:0] n152;
wire      [7:0] n153;
wire      [7:0] n154;
wire      [7:0] n155;
wire      [7:0] n156;
wire      [7:0] n157;
wire      [7:0] n158;
wire     [15:0] n159;
wire     [23:0] n160;
wire     [31:0] n161;
wire     [39:0] n162;
wire     [47:0] n163;
wire     [55:0] n164;
wire     [63:0] n165;
wire     [71:0] n166;
wire      [7:0] n167;
wire      [7:0] n168;
wire      [7:0] n169;
wire      [7:0] n170;
wire      [7:0] n171;
wire      [7:0] n172;
wire      [7:0] n173;
wire      [7:0] n174;
wire      [7:0] n175;
wire     [15:0] n176;
wire     [23:0] n177;
wire     [31:0] n178;
wire     [39:0] n179;
wire     [47:0] n180;
wire     [55:0] n181;
wire     [63:0] n182;
wire     [71:0] n183;
wire      [7:0] n184;
wire      [7:0] n185;
wire      [7:0] n186;
wire      [7:0] n187;
wire      [7:0] n188;
wire      [7:0] n189;
wire      [7:0] n190;
wire      [7:0] n191;
wire      [7:0] n192;
wire     [15:0] n193;
wire     [23:0] n194;
wire     [31:0] n195;
wire     [39:0] n196;
wire     [47:0] n197;
wire     [55:0] n198;
wire     [63:0] n199;
wire     [71:0] n200;
wire    [143:0] n201;
wire    [215:0] n202;
wire    [287:0] n203;
wire    [359:0] n204;
wire    [431:0] n205;
wire    [503:0] n206;
wire    [575:0] n207;
wire    [647:0] n208;
wire    [647:0] n209;
wire    [647:0] n210;
wire      [7:0] n211;
wire      [7:0] n212;
wire      [7:0] n213;
wire      [7:0] n214;
wire      [7:0] n215;
wire      [7:0] n216;
wire            n217;
wire            n218;
wire            n219;
wire            n220;
wire            n221;
wire            n222;
wire            n223;
wire            n224;
wire            n225;
wire            n226;
wire            n227;
wire      [9:0] n228;
wire            n229;
wire            n230;
wire            n231;
wire            n232;
wire            n233;
wire            n234;
wire            n235;
wire            n236;
wire            n237;
wire            n238;
wire            n239;
wire            n240;
wire      [7:0] n241;
wire      [7:0] n242;
wire      [7:0] n243;
wire      [7:0] n244;
wire      [7:0] n245;
wire      [7:0] n246;
wire      [7:0] n247;
wire    [647:0] n248;
wire    [647:0] n249;
wire    [647:0] n250;
wire            n251;
wire            n252;
wire            n253;
wire     [71:0] n254;
wire     [71:0] n255;
wire     [71:0] n256;
wire     [71:0] n257;
wire     [71:0] n258;
wire     [71:0] n259;
wire     [71:0] n260;
wire     [71:0] n261;
wire     [71:0] n262;
wire     [71:0] n263;
wire     [71:0] n264;
wire     [71:0] n265;
wire     [71:0] n266;
wire     [71:0] n267;
wire     [71:0] n268;
wire     [71:0] n269;
wire     [71:0] n270;
wire     [71:0] n271;
wire     [71:0] n272;
wire     [71:0] n273;
wire     [71:0] n274;
wire     [71:0] n275;
wire     [71:0] n276;
wire     [71:0] n277;
wire     [71:0] n278;
wire     [71:0] n279;
wire     [71:0] n280;
wire     [71:0] n281;
wire     [71:0] n282;
wire     [71:0] n283;
wire     [71:0] n284;
wire     [71:0] n285;
wire     [71:0] n286;
wire     [71:0] n287;
wire     [71:0] n288;
wire     [71:0] n289;
wire     [71:0] n290;
wire     [71:0] n291;
wire     [71:0] n292;
wire     [71:0] n293;
wire            n294;
wire      [8:0] n295;
wire      [7:0] n296;
wire            n297;
wire      [7:0] n298;
wire            n299;
wire      [7:0] n300;
wire            n301;
wire      [7:0] n302;
wire            n303;
wire      [7:0] n304;
wire            n305;
wire      [7:0] n306;
wire            n307;
wire      [7:0] n308;
wire      [7:0] n309;
wire      [7:0] n310;
wire      [7:0] n311;
wire      [7:0] n312;
wire      [7:0] n313;
wire      [7:0] n314;
wire      [7:0] n315;
wire      [7:0] n316;
wire      [7:0] n317;
wire      [7:0] n318;
wire      [7:0] n319;
wire      [7:0] n320;
wire      [7:0] n321;
wire      [7:0] n322;
wire      [7:0] n323;
wire      [7:0] n324;
wire      [7:0] n325;
wire      [7:0] n326;
wire      [7:0] n327;
wire      [7:0] n328;
wire      [7:0] n329;
wire      [7:0] n330;
wire      [7:0] n331;
wire      [7:0] n332;
wire      [7:0] n333;
wire      [7:0] n334;
wire      [7:0] n335;
wire      [7:0] n336;
wire      [7:0] n337;
wire      [7:0] n338;
wire      [7:0] n339;
wire      [7:0] n340;
wire      [7:0] n341;
wire      [7:0] n342;
wire      [7:0] n343;
wire      [7:0] n344;
wire      [7:0] n345;
wire      [7:0] n346;
wire      [7:0] n347;
wire      [7:0] n348;
wire      [7:0] n349;
wire      [7:0] n350;
wire      [7:0] n351;
wire      [7:0] n352;
wire      [7:0] n353;
wire      [7:0] n354;
wire      [7:0] n355;
wire      [7:0] n356;
wire      [7:0] n357;
wire      [7:0] n358;
wire      [7:0] n359;
wire      [7:0] n360;
wire      [7:0] n361;
wire      [7:0] n362;
wire      [7:0] n363;
wire      [7:0] n364;
wire      [7:0] n365;
wire     [15:0] n366;
wire     [23:0] n367;
wire     [31:0] n368;
wire     [39:0] n369;
wire     [47:0] n370;
wire     [55:0] n371;
wire     [63:0] n372;
wire     [71:0] n373;
wire     [71:0] n374;
wire     [71:0] n375;
wire     [71:0] n376;
wire     [71:0] n377;
wire     [71:0] n378;
wire      [8:0] RAM_0_addr0;
wire      [7:0] RAM_0_data0;
wire            n379;
wire            n380;
wire            n381;
wire            n382;
wire            n383;
wire            n384;
wire            n385;
wire            n386;
wire            n387;
wire            n388;
wire            n389;
wire            n390;
wire            n391;
wire      [8:0] RAM_1_addr0;
wire      [7:0] RAM_1_data0;
wire            n392;
wire            n393;
wire            n394;
wire      [8:0] RAM_2_addr0;
wire      [7:0] RAM_2_data0;
wire            n395;
wire            n396;
wire            n397;
wire      [8:0] RAM_3_addr0;
wire      [7:0] RAM_3_data0;
wire            n398;
wire            n399;
wire            n400;
wire      [8:0] RAM_4_addr0;
wire      [7:0] RAM_4_data0;
wire            n401;
wire            n402;
wire            n403;
wire      [8:0] RAM_5_addr0;
wire      [7:0] RAM_5_data0;
wire            n404;
wire            n405;
wire            n406;
wire      [8:0] RAM_6_addr0;
wire      [7:0] RAM_6_data0;
wire            n407;
wire            n408;
wire            n409;
wire      [8:0] RAM_7_addr0;
wire      [7:0] RAM_7_data0;
wire            n410;
wire            n411;
wire            n412;
reg      [7:0] RAM_0[511:0];
reg      [7:0] RAM_1[511:0];
reg      [7:0] RAM_2[511:0];
reg      [7:0] RAM_3[511:0];
reg      [7:0] RAM_4[511:0];
reg      [7:0] RAM_5[511:0];
reg      [7:0] RAM_6[511:0];
reg      [7:0] RAM_7[511:0];
wire clk;
wire rst;
wire step;
assign n0 =  ( arg_1_TREADY ) == ( 1'd0 )  ;
assign n1 =  ( arg_0_TVALID ) == ( 1'd0 )  ;
assign n2 =  ( n0 ) & ( n1 )  ;
assign n3 =  ( arg_0_TREADY ) == ( 1'd0 )  ;
assign n4 =  ( n2 ) & ( n3 )  ;
assign n5 =  ( st_ready ) == ( 1'd0 )  ;
assign n6 =  ( n4 ) & ( n5 )  ;
assign n7 =  ( n0 ) & ( n3 )  ;
assign n8 =  ( st_ready ) == ( 1'd1 )  ;
assign n9 =  ( n7 ) & ( n8 )  ;
assign n10 =  ( RAM_x ) == ( 9'd0 )  ;
assign n11 =  ( n9 ) & ( n10 )  ;
assign n12 =  ( RAM_y ) == ( 10'd0 )  ;
assign n13 =  ( n11 ) & ( n12 )  ;
assign n14 =  ( n10 ) & ( n12 )  ;
assign n15 = ~ ( n14 ) ;
assign n16 =  ( n9 ) & ( n15 )  ;
assign n17 =  ( RAM_x ) == ( 9'd488 )  ;
assign n18 =  ( RAM_w ) == ( 3'd7 )  ;
assign n19 =  ( RAM_w ) + ( 3'd1 )  ;
assign n20 =  ( n18 ) ? ( 3'd0 ) : ( n19 ) ;
assign n21 =  ( n17 ) ? ( n20 ) : ( RAM_w ) ;
assign n22 =  ( arg_1_TVALID ) == ( 1'd1 )  ;
assign n23 =  ( arg_1_TREADY ) == ( 1'd1 )  ;
assign n24 =  ( n22 ) & ( n23 )  ;
assign n25 =  ( n24 ) & ( n1 )  ;
assign n26 =  ( n25 ) & ( n3 )  ;
assign n27 =  ( n26 ) ? ( RAM_w ) : ( RAM_w ) ;
assign n28 =  ( n16 ) ? ( n21 ) : ( n27 ) ;
assign n29 =  ( n13 ) ? ( RAM_w ) : ( n28 ) ;
assign n30 =  ( n6 ) ? ( RAM_w ) : ( n29 ) ;
assign n31 =  ( RAM_x ) + ( 9'd1 )  ;
assign n32 =  ( n17 ) ? ( 9'd1 ) : ( n31 ) ;
assign n33 =  ( n26 ) ? ( RAM_x ) : ( RAM_x ) ;
assign n34 =  ( n16 ) ? ( n32 ) : ( n33 ) ;
assign n35 =  ( n13 ) ? ( 9'd1 ) : ( n34 ) ;
assign n36 =  ( n6 ) ? ( RAM_x ) : ( n35 ) ;
assign n37 =  ( RAM_y ) == ( 10'd648 )  ;
assign n38 =  ( RAM_y ) + ( 10'd1 )  ;
assign n39 =  ( n37 ) ? ( 10'd0 ) : ( n38 ) ;
assign n40 =  ( n17 ) ? ( n39 ) : ( RAM_y ) ;
assign n41 =  ( n26 ) ? ( RAM_y ) : ( RAM_y ) ;
assign n42 =  ( n16 ) ? ( n40 ) : ( n41 ) ;
assign n43 =  ( n13 ) ? ( RAM_y ) : ( n42 ) ;
assign n44 =  ( n6 ) ? ( RAM_y ) : ( n43 ) ;
assign n45 =  ( RAM_x ) == ( 9'd1 )  ;
assign n46 =  ( n45 ) & ( n37 )  ;
assign n47 =  ( RAM_x ) > ( 9'd8 )  ;
assign n48 = stencil_8[71:64] ;
assign n49 = stencil_7[71:64] ;
assign n50 = stencil_6[71:64] ;
assign n51 = stencil_5[71:64] ;
assign n52 = stencil_4[71:64] ;
assign n53 = stencil_3[71:64] ;
assign n54 = stencil_2[71:64] ;
assign n55 = stencil_1[71:64] ;
assign n56 = stencil_0[71:64] ;
assign n57 =  { ( n55 ) , ( n56 ) }  ;
assign n58 =  { ( n54 ) , ( n57 ) }  ;
assign n59 =  { ( n53 ) , ( n58 ) }  ;
assign n60 =  { ( n52 ) , ( n59 ) }  ;
assign n61 =  { ( n51 ) , ( n60 ) }  ;
assign n62 =  { ( n50 ) , ( n61 ) }  ;
assign n63 =  { ( n49 ) , ( n62 ) }  ;
assign n64 =  { ( n48 ) , ( n63 ) }  ;
assign n65 = stencil_8[63:56] ;
assign n66 = stencil_7[63:56] ;
assign n67 = stencil_6[63:56] ;
assign n68 = stencil_5[63:56] ;
assign n69 = stencil_4[63:56] ;
assign n70 = stencil_3[63:56] ;
assign n71 = stencil_2[63:56] ;
assign n72 = stencil_1[63:56] ;
assign n73 = stencil_0[63:56] ;
assign n74 =  { ( n72 ) , ( n73 ) }  ;
assign n75 =  { ( n71 ) , ( n74 ) }  ;
assign n76 =  { ( n70 ) , ( n75 ) }  ;
assign n77 =  { ( n69 ) , ( n76 ) }  ;
assign n78 =  { ( n68 ) , ( n77 ) }  ;
assign n79 =  { ( n67 ) , ( n78 ) }  ;
assign n80 =  { ( n66 ) , ( n79 ) }  ;
assign n81 =  { ( n65 ) , ( n80 ) }  ;
assign n82 = stencil_8[55:48] ;
assign n83 = stencil_7[55:48] ;
assign n84 = stencil_6[55:48] ;
assign n85 = stencil_5[55:48] ;
assign n86 = stencil_4[55:48] ;
assign n87 = stencil_3[55:48] ;
assign n88 = stencil_2[55:48] ;
assign n89 = stencil_1[55:48] ;
assign n90 = stencil_0[55:48] ;
assign n91 =  { ( n89 ) , ( n90 ) }  ;
assign n92 =  { ( n88 ) , ( n91 ) }  ;
assign n93 =  { ( n87 ) , ( n92 ) }  ;
assign n94 =  { ( n86 ) , ( n93 ) }  ;
assign n95 =  { ( n85 ) , ( n94 ) }  ;
assign n96 =  { ( n84 ) , ( n95 ) }  ;
assign n97 =  { ( n83 ) , ( n96 ) }  ;
assign n98 =  { ( n82 ) , ( n97 ) }  ;
assign n99 = stencil_8[47:40] ;
assign n100 = stencil_7[47:40] ;
assign n101 = stencil_6[47:40] ;
assign n102 = stencil_5[47:40] ;
assign n103 = stencil_4[47:40] ;
assign n104 = stencil_3[47:40] ;
assign n105 = stencil_2[47:40] ;
assign n106 = stencil_1[47:40] ;
assign n107 = stencil_0[47:40] ;
assign n108 =  { ( n106 ) , ( n107 ) }  ;
assign n109 =  { ( n105 ) , ( n108 ) }  ;
assign n110 =  { ( n104 ) , ( n109 ) }  ;
assign n111 =  { ( n103 ) , ( n110 ) }  ;
assign n112 =  { ( n102 ) , ( n111 ) }  ;
assign n113 =  { ( n101 ) , ( n112 ) }  ;
assign n114 =  { ( n100 ) , ( n113 ) }  ;
assign n115 =  { ( n99 ) , ( n114 ) }  ;
assign n116 = stencil_8[39:32] ;
assign n117 = stencil_7[39:32] ;
assign n118 = stencil_6[39:32] ;
assign n119 = stencil_5[39:32] ;
assign n120 = stencil_4[39:32] ;
assign n121 = stencil_3[39:32] ;
assign n122 = stencil_2[39:32] ;
assign n123 = stencil_1[39:32] ;
assign n124 = stencil_0[39:32] ;
assign n125 =  { ( n123 ) , ( n124 ) }  ;
assign n126 =  { ( n122 ) , ( n125 ) }  ;
assign n127 =  { ( n121 ) , ( n126 ) }  ;
assign n128 =  { ( n120 ) , ( n127 ) }  ;
assign n129 =  { ( n119 ) , ( n128 ) }  ;
assign n130 =  { ( n118 ) , ( n129 ) }  ;
assign n131 =  { ( n117 ) , ( n130 ) }  ;
assign n132 =  { ( n116 ) , ( n131 ) }  ;
assign n133 = stencil_8[31:24] ;
assign n134 = stencil_7[31:24] ;
assign n135 = stencil_6[31:24] ;
assign n136 = stencil_5[31:24] ;
assign n137 = stencil_4[31:24] ;
assign n138 = stencil_3[31:24] ;
assign n139 = stencil_2[31:24] ;
assign n140 = stencil_1[31:24] ;
assign n141 = stencil_0[31:24] ;
assign n142 =  { ( n140 ) , ( n141 ) }  ;
assign n143 =  { ( n139 ) , ( n142 ) }  ;
assign n144 =  { ( n138 ) , ( n143 ) }  ;
assign n145 =  { ( n137 ) , ( n144 ) }  ;
assign n146 =  { ( n136 ) , ( n145 ) }  ;
assign n147 =  { ( n135 ) , ( n146 ) }  ;
assign n148 =  { ( n134 ) , ( n147 ) }  ;
assign n149 =  { ( n133 ) , ( n148 ) }  ;
assign n150 = stencil_8[23:16] ;
assign n151 = stencil_7[23:16] ;
assign n152 = stencil_6[23:16] ;
assign n153 = stencil_5[23:16] ;
assign n154 = stencil_4[23:16] ;
assign n155 = stencil_3[23:16] ;
assign n156 = stencil_2[23:16] ;
assign n157 = stencil_1[23:16] ;
assign n158 = stencil_0[23:16] ;
assign n159 =  { ( n157 ) , ( n158 ) }  ;
assign n160 =  { ( n156 ) , ( n159 ) }  ;
assign n161 =  { ( n155 ) , ( n160 ) }  ;
assign n162 =  { ( n154 ) , ( n161 ) }  ;
assign n163 =  { ( n153 ) , ( n162 ) }  ;
assign n164 =  { ( n152 ) , ( n163 ) }  ;
assign n165 =  { ( n151 ) , ( n164 ) }  ;
assign n166 =  { ( n150 ) , ( n165 ) }  ;
assign n167 = stencil_8[15:8] ;
assign n168 = stencil_7[15:8] ;
assign n169 = stencil_6[15:8] ;
assign n170 = stencil_5[15:8] ;
assign n171 = stencil_4[15:8] ;
assign n172 = stencil_3[15:8] ;
assign n173 = stencil_2[15:8] ;
assign n174 = stencil_1[15:8] ;
assign n175 = stencil_0[15:8] ;
assign n176 =  { ( n174 ) , ( n175 ) }  ;
assign n177 =  { ( n173 ) , ( n176 ) }  ;
assign n178 =  { ( n172 ) , ( n177 ) }  ;
assign n179 =  { ( n171 ) , ( n178 ) }  ;
assign n180 =  { ( n170 ) , ( n179 ) }  ;
assign n181 =  { ( n169 ) , ( n180 ) }  ;
assign n182 =  { ( n168 ) , ( n181 ) }  ;
assign n183 =  { ( n167 ) , ( n182 ) }  ;
assign n184 = stencil_8[7:0] ;
assign n185 = stencil_7[7:0] ;
assign n186 = stencil_6[7:0] ;
assign n187 = stencil_5[7:0] ;
assign n188 = stencil_4[7:0] ;
assign n189 = stencil_3[7:0] ;
assign n190 = stencil_2[7:0] ;
assign n191 = stencil_1[7:0] ;
assign n192 = stencil_0[7:0] ;
assign n193 =  { ( n191 ) , ( n192 ) }  ;
assign n194 =  { ( n190 ) , ( n193 ) }  ;
assign n195 =  { ( n189 ) , ( n194 ) }  ;
assign n196 =  { ( n188 ) , ( n195 ) }  ;
assign n197 =  { ( n187 ) , ( n196 ) }  ;
assign n198 =  { ( n186 ) , ( n197 ) }  ;
assign n199 =  { ( n185 ) , ( n198 ) }  ;
assign n200 =  { ( n184 ) , ( n199 ) }  ;
assign n201 =  { ( n183 ) , ( n200 ) }  ;
assign n202 =  { ( n166 ) , ( n201 ) }  ;
assign n203 =  { ( n149 ) , ( n202 ) }  ;
assign n204 =  { ( n132 ) , ( n203 ) }  ;
assign n205 =  { ( n115 ) , ( n204 ) }  ;
assign n206 =  { ( n98 ) , ( n205 ) }  ;
assign n207 =  { ( n81 ) , ( n206 ) }  ;
assign n208 =  { ( n64 ) , ( n207 ) }  ;
assign n209 =  ( n47 ) ? ( n208 ) : ( proc_in ) ;
assign n210 =  ( n46 ) ? ( proc_in ) : ( n209 ) ;
assign n211 = gb_fun(n210) ;
assign n212 =  ( n46 ) ? ( arg_0_TDATA ) : ( n211 ) ;
assign n213 =  ( n26 ) ? ( arg_0_TDATA ) : ( arg_0_TDATA ) ;
assign n214 =  ( n16 ) ? ( arg_0_TDATA ) : ( n213 ) ;
assign n215 =  ( n13 ) ? ( arg_0_TDATA ) : ( n214 ) ;
assign n216 =  ( n6 ) ? ( n212 ) : ( n215 ) ;
assign n217 =  ( RAM_y ) >= ( 10'd8 )  ;
assign n218 =  ( n47 ) & ( n217 )  ;
assign n219 =  ( RAM_y ) > ( 10'd8 )  ;
assign n220 =  ( n45 ) & ( n219 )  ;
assign n221 =  ( n218 ) | ( n220 )  ;
assign n222 =  ( n221 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n223 =  ( n46 ) ? ( arg_0_TVALID ) : ( n222 ) ;
assign n224 =  ( n26 ) ? ( 1'd0 ) : ( arg_0_TVALID ) ;
assign n225 =  ( n16 ) ? ( arg_0_TVALID ) : ( n224 ) ;
assign n226 =  ( n13 ) ? ( 1'd0 ) : ( n225 ) ;
assign n227 =  ( n6 ) ? ( n223 ) : ( n226 ) ;
assign n228 =  ( 10'd648 ) - ( 10'd1 )  ;
assign n229 =  ( RAM_y ) == ( n228 )  ;
assign n230 =  ( n17 ) & ( n229 )  ;
assign n231 =  ( n230 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n232 =  ( RAM_y ) < ( 10'd8 )  ;
assign n233 =  ( RAM_y ) == ( 10'd8 )  ;
assign n234 =  ( n233 ) & ( n45 )  ;
assign n235 =  ( n232 ) | ( n234 )  ;
assign n236 =  ( n235 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n237 =  ( n26 ) ? ( 1'd0 ) : ( arg_1_TREADY ) ;
assign n238 =  ( n16 ) ? ( n236 ) : ( n237 ) ;
assign n239 =  ( n13 ) ? ( 1'd1 ) : ( n238 ) ;
assign n240 =  ( n6 ) ? ( n231 ) : ( n239 ) ;
assign n241 =  ( n26 ) ? ( arg_1_TDATA ) : ( cur_pix ) ;
assign n242 =  ( n16 ) ? ( cur_pix ) : ( n241 ) ;
assign n243 =  ( n13 ) ? ( cur_pix ) : ( n242 ) ;
assign n244 =  ( n6 ) ? ( cur_pix ) : ( n243 ) ;
assign n245 =  ( n16 ) ? ( cur_pix ) : ( pre_pix ) ;
assign n246 =  ( n13 ) ? ( cur_pix ) : ( n245 ) ;
assign n247 =  ( n6 ) ? ( pre_pix ) : ( n246 ) ;
assign n248 =  ( n16 ) ? ( proc_in ) : ( proc_in ) ;
assign n249 =  ( n13 ) ? ( proc_in ) : ( n248 ) ;
assign n250 =  ( n6 ) ? ( n210 ) : ( n249 ) ;
assign n251 =  ( n16 ) ? ( n236 ) : ( st_ready ) ;
assign n252 =  ( n13 ) ? ( 1'd1 ) : ( n251 ) ;
assign n253 =  ( n6 ) ? ( 1'd1 ) : ( n252 ) ;
assign n254 =  ( n232 ) ? ( stencil_0 ) : ( stencil_1 ) ;
assign n255 =  ( n26 ) ? ( stencil_0 ) : ( stencil_0 ) ;
assign n256 =  ( n16 ) ? ( stencil_0 ) : ( n255 ) ;
assign n257 =  ( n13 ) ? ( stencil_0 ) : ( n256 ) ;
assign n258 =  ( n6 ) ? ( n254 ) : ( n257 ) ;
assign n259 =  ( n232 ) ? ( stencil_1 ) : ( stencil_2 ) ;
assign n260 =  ( n26 ) ? ( stencil_1 ) : ( stencil_1 ) ;
assign n261 =  ( n16 ) ? ( stencil_1 ) : ( n260 ) ;
assign n262 =  ( n13 ) ? ( stencil_1 ) : ( n261 ) ;
assign n263 =  ( n6 ) ? ( n259 ) : ( n262 ) ;
assign n264 =  ( n232 ) ? ( stencil_2 ) : ( stencil_3 ) ;
assign n265 =  ( n26 ) ? ( stencil_2 ) : ( stencil_2 ) ;
assign n266 =  ( n16 ) ? ( stencil_2 ) : ( n265 ) ;
assign n267 =  ( n13 ) ? ( stencil_2 ) : ( n266 ) ;
assign n268 =  ( n6 ) ? ( n264 ) : ( n267 ) ;
assign n269 =  ( n232 ) ? ( stencil_3 ) : ( stencil_4 ) ;
assign n270 =  ( n26 ) ? ( stencil_3 ) : ( stencil_3 ) ;
assign n271 =  ( n16 ) ? ( stencil_3 ) : ( n270 ) ;
assign n272 =  ( n13 ) ? ( stencil_3 ) : ( n271 ) ;
assign n273 =  ( n6 ) ? ( n269 ) : ( n272 ) ;
assign n274 =  ( n232 ) ? ( stencil_4 ) : ( stencil_5 ) ;
assign n275 =  ( n26 ) ? ( stencil_4 ) : ( stencil_4 ) ;
assign n276 =  ( n16 ) ? ( stencil_4 ) : ( n275 ) ;
assign n277 =  ( n13 ) ? ( stencil_4 ) : ( n276 ) ;
assign n278 =  ( n6 ) ? ( n274 ) : ( n277 ) ;
assign n279 =  ( n232 ) ? ( stencil_5 ) : ( stencil_6 ) ;
assign n280 =  ( n26 ) ? ( stencil_5 ) : ( stencil_5 ) ;
assign n281 =  ( n16 ) ? ( stencil_5 ) : ( n280 ) ;
assign n282 =  ( n13 ) ? ( stencil_5 ) : ( n281 ) ;
assign n283 =  ( n6 ) ? ( n279 ) : ( n282 ) ;
assign n284 =  ( n232 ) ? ( stencil_6 ) : ( stencil_7 ) ;
assign n285 =  ( n26 ) ? ( stencil_6 ) : ( stencil_6 ) ;
assign n286 =  ( n16 ) ? ( stencil_6 ) : ( n285 ) ;
assign n287 =  ( n13 ) ? ( stencil_6 ) : ( n286 ) ;
assign n288 =  ( n6 ) ? ( n284 ) : ( n287 ) ;
assign n289 =  ( n232 ) ? ( stencil_7 ) : ( stencil_8 ) ;
assign n290 =  ( n26 ) ? ( stencil_7 ) : ( stencil_7 ) ;
assign n291 =  ( n16 ) ? ( stencil_7 ) : ( n290 ) ;
assign n292 =  ( n13 ) ? ( stencil_7 ) : ( n291 ) ;
assign n293 =  ( n6 ) ? ( n289 ) : ( n292 ) ;
assign n294 =  ( RAM_w ) == ( 3'd0 )  ;
assign n295 =  ( RAM_x ) - ( 9'd1 )  ;
assign n296 =  (  RAM_7 [ n295 ] )  ;
assign n297 =  ( RAM_w ) == ( 3'd1 )  ;
assign n298 =  (  RAM_0 [ n295 ] )  ;
assign n299 =  ( RAM_w ) == ( 3'd2 )  ;
assign n300 =  (  RAM_1 [ n295 ] )  ;
assign n301 =  ( RAM_w ) == ( 3'd3 )  ;
assign n302 =  (  RAM_2 [ n295 ] )  ;
assign n303 =  ( RAM_w ) == ( 3'd4 )  ;
assign n304 =  (  RAM_3 [ n295 ] )  ;
assign n305 =  ( RAM_w ) == ( 3'd5 )  ;
assign n306 =  (  RAM_4 [ n295 ] )  ;
assign n307 =  ( RAM_w ) == ( 3'd6 )  ;
assign n308 =  (  RAM_5 [ n295 ] )  ;
assign n309 =  (  RAM_6 [ n295 ] )  ;
assign n310 =  ( n307 ) ? ( n308 ) : ( n309 ) ;
assign n311 =  ( n305 ) ? ( n306 ) : ( n310 ) ;
assign n312 =  ( n303 ) ? ( n304 ) : ( n311 ) ;
assign n313 =  ( n301 ) ? ( n302 ) : ( n312 ) ;
assign n314 =  ( n299 ) ? ( n300 ) : ( n313 ) ;
assign n315 =  ( n297 ) ? ( n298 ) : ( n314 ) ;
assign n316 =  ( n294 ) ? ( n296 ) : ( n315 ) ;
assign n317 =  ( n307 ) ? ( n306 ) : ( n308 ) ;
assign n318 =  ( n305 ) ? ( n304 ) : ( n317 ) ;
assign n319 =  ( n303 ) ? ( n302 ) : ( n318 ) ;
assign n320 =  ( n301 ) ? ( n300 ) : ( n319 ) ;
assign n321 =  ( n299 ) ? ( n298 ) : ( n320 ) ;
assign n322 =  ( n297 ) ? ( n296 ) : ( n321 ) ;
assign n323 =  ( n294 ) ? ( n309 ) : ( n322 ) ;
assign n324 =  ( n307 ) ? ( n304 ) : ( n306 ) ;
assign n325 =  ( n305 ) ? ( n302 ) : ( n324 ) ;
assign n326 =  ( n303 ) ? ( n300 ) : ( n325 ) ;
assign n327 =  ( n301 ) ? ( n298 ) : ( n326 ) ;
assign n328 =  ( n299 ) ? ( n296 ) : ( n327 ) ;
assign n329 =  ( n297 ) ? ( n309 ) : ( n328 ) ;
assign n330 =  ( n294 ) ? ( n308 ) : ( n329 ) ;
assign n331 =  ( n307 ) ? ( n302 ) : ( n304 ) ;
assign n332 =  ( n305 ) ? ( n300 ) : ( n331 ) ;
assign n333 =  ( n303 ) ? ( n298 ) : ( n332 ) ;
assign n334 =  ( n301 ) ? ( n296 ) : ( n333 ) ;
assign n335 =  ( n299 ) ? ( n309 ) : ( n334 ) ;
assign n336 =  ( n297 ) ? ( n308 ) : ( n335 ) ;
assign n337 =  ( n294 ) ? ( n306 ) : ( n336 ) ;
assign n338 =  ( n307 ) ? ( n300 ) : ( n302 ) ;
assign n339 =  ( n305 ) ? ( n298 ) : ( n338 ) ;
assign n340 =  ( n303 ) ? ( n296 ) : ( n339 ) ;
assign n341 =  ( n301 ) ? ( n309 ) : ( n340 ) ;
assign n342 =  ( n299 ) ? ( n308 ) : ( n341 ) ;
assign n343 =  ( n297 ) ? ( n306 ) : ( n342 ) ;
assign n344 =  ( n294 ) ? ( n304 ) : ( n343 ) ;
assign n345 =  ( n307 ) ? ( n298 ) : ( n300 ) ;
assign n346 =  ( n305 ) ? ( n296 ) : ( n345 ) ;
assign n347 =  ( n303 ) ? ( n309 ) : ( n346 ) ;
assign n348 =  ( n301 ) ? ( n308 ) : ( n347 ) ;
assign n349 =  ( n299 ) ? ( n306 ) : ( n348 ) ;
assign n350 =  ( n297 ) ? ( n304 ) : ( n349 ) ;
assign n351 =  ( n294 ) ? ( n302 ) : ( n350 ) ;
assign n352 =  ( n307 ) ? ( n296 ) : ( n298 ) ;
assign n353 =  ( n305 ) ? ( n309 ) : ( n352 ) ;
assign n354 =  ( n303 ) ? ( n308 ) : ( n353 ) ;
assign n355 =  ( n301 ) ? ( n306 ) : ( n354 ) ;
assign n356 =  ( n299 ) ? ( n304 ) : ( n355 ) ;
assign n357 =  ( n297 ) ? ( n302 ) : ( n356 ) ;
assign n358 =  ( n294 ) ? ( n300 ) : ( n357 ) ;
assign n359 =  ( n307 ) ? ( n309 ) : ( n296 ) ;
assign n360 =  ( n305 ) ? ( n308 ) : ( n359 ) ;
assign n361 =  ( n303 ) ? ( n306 ) : ( n360 ) ;
assign n362 =  ( n301 ) ? ( n304 ) : ( n361 ) ;
assign n363 =  ( n299 ) ? ( n302 ) : ( n362 ) ;
assign n364 =  ( n297 ) ? ( n300 ) : ( n363 ) ;
assign n365 =  ( n294 ) ? ( n298 ) : ( n364 ) ;
assign n366 =  { ( n358 ) , ( n365 ) }  ;
assign n367 =  { ( n351 ) , ( n366 ) }  ;
assign n368 =  { ( n344 ) , ( n367 ) }  ;
assign n369 =  { ( n337 ) , ( n368 ) }  ;
assign n370 =  { ( n330 ) , ( n369 ) }  ;
assign n371 =  { ( n323 ) , ( n370 ) }  ;
assign n372 =  { ( n316 ) , ( n371 ) }  ;
assign n373 =  { ( pre_pix ) , ( n372 ) }  ;
assign n374 =  ( n232 ) ? ( stencil_8 ) : ( n373 ) ;
assign n375 =  ( n26 ) ? ( stencil_8 ) : ( stencil_8 ) ;
assign n376 =  ( n16 ) ? ( n374 ) : ( n375 ) ;
assign n377 =  ( n13 ) ? ( stencil_8 ) : ( n376 ) ;
assign n378 =  ( n6 ) ? ( stencil_8 ) : ( n377 ) ;
assign n379 = ~ ( n6 ) ;
assign n380 = ~ ( n13 ) ;
assign n381 =  ( n379 ) & ( n380 )  ;
assign n382 = ~ ( n16 ) ;
assign n383 =  ( n381 ) & ( n382 )  ;
assign n384 = ~ ( n26 ) ;
assign n385 =  ( n383 ) & ( n384 )  ;
assign n386 =  ( n383 ) & ( n26 )  ;
assign n387 =  ( n381 ) & ( n16 )  ;
assign n388 = ~ ( n294 ) ;
assign n389 =  ( n387 ) & ( n388 )  ;
assign n390 =  ( n387 ) & ( n294 )  ;
assign n391 =  ( n379 ) & ( n13 )  ;
assign RAM_0_addr0 = n390 ? (n295) : (0);
assign RAM_0_data0 = n390 ? (pre_pix) : (RAM_0[0]);
assign n392 = ~ ( n297 ) ;
assign n393 =  ( n387 ) & ( n392 )  ;
assign n394 =  ( n387 ) & ( n297 )  ;
assign RAM_1_addr0 = n394 ? (n295) : (0);
assign RAM_1_data0 = n394 ? (pre_pix) : (RAM_1[0]);
assign n395 = ~ ( n299 ) ;
assign n396 =  ( n387 ) & ( n395 )  ;
assign n397 =  ( n387 ) & ( n299 )  ;
assign RAM_2_addr0 = n397 ? (n295) : (0);
assign RAM_2_data0 = n397 ? (pre_pix) : (RAM_2[0]);
assign n398 = ~ ( n301 ) ;
assign n399 =  ( n387 ) & ( n398 )  ;
assign n400 =  ( n387 ) & ( n301 )  ;
assign RAM_3_addr0 = n400 ? (n295) : (0);
assign RAM_3_data0 = n400 ? (pre_pix) : (RAM_3[0]);
assign n401 = ~ ( n303 ) ;
assign n402 =  ( n387 ) & ( n401 )  ;
assign n403 =  ( n387 ) & ( n303 )  ;
assign RAM_4_addr0 = n403 ? (n295) : (0);
assign RAM_4_data0 = n403 ? (pre_pix) : (RAM_4[0]);
assign n404 = ~ ( n305 ) ;
assign n405 =  ( n387 ) & ( n404 )  ;
assign n406 =  ( n387 ) & ( n305 )  ;
assign RAM_5_addr0 = n406 ? (n295) : (0);
assign RAM_5_data0 = n406 ? (pre_pix) : (RAM_5[0]);
assign n407 = ~ ( n307 ) ;
assign n408 =  ( n387 ) & ( n407 )  ;
assign n409 =  ( n387 ) & ( n307 )  ;
assign RAM_6_addr0 = n409 ? (n295) : (0);
assign RAM_6_data0 = n409 ? (pre_pix) : (RAM_6[0]);
assign n410 = ~ ( n18 ) ;
assign n411 =  ( n387 ) & ( n410 )  ;
assign n412 =  ( n387 ) & ( n18 )  ;
assign RAM_7_addr0 = n412 ? (n295) : (0);
assign RAM_7_data0 = n412 ? (pre_pix) : (RAM_7[0]);
function [7:0] gb_fun ;
input [647:0] arg0;
    begin
//TODO: Add the specific function HERE.    end
endfunction

always @(posedge clk) begin
   if(rst) begin
       RAM_w <= RAM_w;
       RAM_x <= RAM_x;
       RAM_y <= RAM_y;
       arg_0_TDATA <= arg_0_TDATA;
       arg_0_TVALID <= arg_0_TVALID;
       arg_1_TREADY <= arg_1_TREADY;
       cur_pix <= cur_pix;
       pre_pix <= pre_pix;
       proc_in <= proc_in;
       st_ready <= st_ready;
       stencil_0 <= stencil_0;
       stencil_1 <= stencil_1;
       stencil_2 <= stencil_2;
       stencil_3 <= stencil_3;
       stencil_4 <= stencil_4;
       stencil_5 <= stencil_5;
       stencil_6 <= stencil_6;
       stencil_7 <= stencil_7;
       stencil_8 <= stencil_8;
   end
   else if(step) begin
       RAM_w <= n30;
       RAM_x <= n36;
       RAM_y <= n44;
       arg_0_TDATA <= n216;
       arg_0_TVALID <= n227;
       arg_1_TREADY <= n240;
       cur_pix <= n244;
       pre_pix <= n247;
       proc_in <= n250;
       st_ready <= n253;
       stencil_0 <= n258;
       stencil_1 <= n263;
       stencil_2 <= n268;
       stencil_3 <= n273;
       stencil_4 <= n278;
       stencil_5 <= n283;
       stencil_6 <= n288;
       stencil_7 <= n293;
       stencil_8 <= n378;
       RAM_0 [ RAM_0_addr0 ] <= RAM_0_data0;
       RAM_1 [ RAM_1_addr0 ] <= RAM_1_data0;
       RAM_2 [ RAM_2_addr0 ] <= RAM_2_data0;
       RAM_3 [ RAM_3_addr0 ] <= RAM_3_data0;
       RAM_4 [ RAM_4_addr0 ] <= RAM_4_data0;
       RAM_5 [ RAM_5_addr0 ] <= RAM_5_data0;
       RAM_6 [ RAM_6_addr0 ] <= RAM_6_data0;
       RAM_7 [ RAM_7_addr0 ] <= RAM_7_data0;
   end
end
endmodule
