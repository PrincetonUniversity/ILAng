module A(
    input clk,
    input rst, output r);

`include "m2.v"    
    
endmodule

