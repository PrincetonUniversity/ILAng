module GB(
arg_0_TREADY,
arg_1_TDATA,
arg_1_TVALID,
LB1D_buff,
LB1D_p_cnt,
LB2D_proc_w,
LB2D_proc_x,
LB2D_proc_y,
LB2D_shift_0,
LB2D_shift_1,
LB2D_shift_2,
LB2D_shift_3,
LB2D_shift_4,
LB2D_shift_5,
LB2D_shift_6,
LB2D_shift_7,
LB2D_shift_x,
LB2D_shift_y,
arg_0_TDATA,
arg_0_TVALID,
arg_1_TREADY,
gb_exit_it_1,
gb_exit_it_2,
gb_exit_it_3,
gb_exit_it_4,
gb_exit_it_5,
gb_exit_it_6,
gb_exit_it_7,
gb_exit_it_8,
gb_p_cnt,
gb_pp_it_1,
gb_pp_it_2,
gb_pp_it_3,
gb_pp_it_4,
gb_pp_it_5,
gb_pp_it_6,
gb_pp_it_7,
gb_pp_it_8,
gb_pp_it_9,
in_stream_buff_0,
in_stream_buff_1,
in_stream_empty,
in_stream_full,
slice_stream_buff_0,
slice_stream_buff_1,
slice_stream_empty,
slice_stream_full,
stencil_stream_buff_0,
stencil_stream_buff_1,
stencil_stream_empty,
stencil_stream_full,
clk,rst,
step
);
input            arg_0_TREADY;
input      [7:0] arg_1_TDATA;
input            arg_1_TVALID;
input clk;
input rst;
input step;
output      [7:0] LB1D_buff;
output     [18:0] LB1D_p_cnt;
output     [63:0] LB2D_proc_w;
output      [8:0] LB2D_proc_x;
output      [9:0] LB2D_proc_y;
output     [71:0] LB2D_shift_0;
output     [71:0] LB2D_shift_1;
output     [71:0] LB2D_shift_2;
output     [71:0] LB2D_shift_3;
output     [71:0] LB2D_shift_4;
output     [71:0] LB2D_shift_5;
output     [71:0] LB2D_shift_6;
output     [71:0] LB2D_shift_7;
output      [8:0] LB2D_shift_x;
output      [9:0] LB2D_shift_y;
output      [7:0] arg_0_TDATA;
output            arg_0_TVALID;
output            arg_1_TREADY;
output            gb_exit_it_1;
output            gb_exit_it_2;
output            gb_exit_it_3;
output            gb_exit_it_4;
output            gb_exit_it_5;
output            gb_exit_it_6;
output            gb_exit_it_7;
output            gb_exit_it_8;
output     [18:0] gb_p_cnt;
output            gb_pp_it_1;
output            gb_pp_it_2;
output            gb_pp_it_3;
output            gb_pp_it_4;
output            gb_pp_it_5;
output            gb_pp_it_6;
output            gb_pp_it_7;
output            gb_pp_it_8;
output            gb_pp_it_9;
output      [7:0] in_stream_buff_0;
output      [7:0] in_stream_buff_1;
output            in_stream_empty;
output            in_stream_full;
output     [71:0] slice_stream_buff_0;
output     [71:0] slice_stream_buff_1;
output            slice_stream_empty;
output            slice_stream_full;
output    [647:0] stencil_stream_buff_0;
output    [647:0] stencil_stream_buff_1;
output            stencil_stream_empty;
output            stencil_stream_full;
reg      [7:0] LB1D_buff;
reg     [18:0] LB1D_p_cnt;
reg     [63:0] LB2D_proc_w;
reg      [8:0] LB2D_proc_x;
reg      [9:0] LB2D_proc_y;
reg     [71:0] LB2D_shift_0;
reg     [71:0] LB2D_shift_1;
reg     [71:0] LB2D_shift_2;
reg     [71:0] LB2D_shift_3;
reg     [71:0] LB2D_shift_4;
reg     [71:0] LB2D_shift_5;
reg     [71:0] LB2D_shift_6;
reg     [71:0] LB2D_shift_7;
reg      [8:0] LB2D_shift_x;
reg      [9:0] LB2D_shift_y;
reg      [7:0] arg_0_TDATA;
reg            arg_0_TVALID;
reg            arg_1_TREADY;
reg            gb_exit_it_1;
reg            gb_exit_it_2;
reg            gb_exit_it_3;
reg            gb_exit_it_4;
reg            gb_exit_it_5;
reg            gb_exit_it_6;
reg            gb_exit_it_7;
reg            gb_exit_it_8;
reg     [18:0] gb_p_cnt;
reg            gb_pp_it_1;
reg            gb_pp_it_2;
reg            gb_pp_it_3;
reg            gb_pp_it_4;
reg            gb_pp_it_5;
reg            gb_pp_it_6;
reg            gb_pp_it_7;
reg            gb_pp_it_8;
reg            gb_pp_it_9;
reg      [7:0] in_stream_buff_0;
reg      [7:0] in_stream_buff_1;
reg            in_stream_empty;
reg            in_stream_full;
reg     [71:0] slice_stream_buff_0;
reg     [71:0] slice_stream_buff_1;
reg            slice_stream_empty;
reg            slice_stream_full;
reg    [647:0] stencil_stream_buff_0;
reg    [647:0] stencil_stream_buff_1;
reg            stencil_stream_empty;
reg            stencil_stream_full;
wire            arg_0_TREADY;
wire      [7:0] arg_1_TDATA;
wire            arg_1_TVALID;
wire            n0;
wire            n1;
wire            n2;
wire            n3;
wire            n4;
wire            n5;
wire            n6;
wire            n7;
wire            n8;
wire            n9;
wire            n10;
wire            n11;
wire            n12;
wire            n13;
wire            n14;
wire            n15;
wire            n16;
wire            n17;
wire            n18;
wire            n19;
wire            n20;
wire            n21;
wire            n22;
wire            n23;
wire            n24;
wire            n25;
wire            n26;
wire            n27;
wire            n28;
wire            n29;
wire            n30;
wire            n31;
wire            n32;
wire            n33;
wire            n34;
wire            n35;
wire      [7:0] n36;
wire      [7:0] n37;
wire      [7:0] n38;
wire      [7:0] n39;
wire      [7:0] n40;
wire      [7:0] n41;
wire     [18:0] n42;
wire     [18:0] n43;
wire     [18:0] n44;
wire     [18:0] n45;
wire     [18:0] n46;
wire     [18:0] n47;
wire     [18:0] n48;
wire            n49;
wire            n50;
wire     [63:0] n51;
wire     [63:0] n52;
wire     [63:0] n53;
wire     [63:0] n54;
wire     [63:0] n55;
wire     [63:0] n56;
wire     [63:0] n57;
wire     [63:0] n58;
wire     [63:0] n59;
wire            n60;
wire            n61;
wire            n62;
wire      [8:0] n63;
wire      [8:0] n64;
wire      [8:0] n65;
wire      [8:0] n66;
wire      [8:0] n67;
wire      [8:0] n68;
wire      [8:0] n69;
wire      [8:0] n70;
wire            n71;
wire      [9:0] n72;
wire      [9:0] n73;
wire      [9:0] n74;
wire      [9:0] n75;
wire      [9:0] n76;
wire      [9:0] n77;
wire      [9:0] n78;
wire            n79;
wire     [71:0] n80;
wire     [71:0] n81;
wire     [71:0] n82;
wire     [71:0] n83;
wire     [71:0] n84;
wire     [71:0] n85;
wire     [71:0] n86;
wire     [71:0] n87;
wire     [71:0] n88;
wire     [71:0] n89;
wire     [71:0] n90;
wire     [71:0] n91;
wire     [71:0] n92;
wire     [71:0] n93;
wire     [71:0] n94;
wire     [71:0] n95;
wire     [71:0] n96;
wire     [71:0] n97;
wire     [71:0] n98;
wire     [71:0] n99;
wire     [71:0] n100;
wire     [71:0] n101;
wire     [71:0] n102;
wire     [71:0] n103;
wire     [71:0] n104;
wire     [71:0] n105;
wire     [71:0] n106;
wire     [71:0] n107;
wire     [71:0] n108;
wire     [71:0] n109;
wire     [71:0] n110;
wire     [71:0] n111;
wire     [71:0] n112;
wire     [71:0] n113;
wire     [71:0] n114;
wire     [71:0] n115;
wire     [71:0] n116;
wire     [71:0] n117;
wire     [71:0] n118;
wire     [71:0] n119;
wire     [71:0] n120;
wire     [71:0] n121;
wire     [71:0] n122;
wire     [71:0] n123;
wire     [71:0] n124;
wire     [71:0] n125;
wire     [71:0] n126;
wire     [71:0] n127;
wire     [71:0] n128;
wire            n129;
wire      [8:0] n130;
wire      [8:0] n131;
wire      [8:0] n132;
wire      [8:0] n133;
wire      [8:0] n134;
wire      [8:0] n135;
wire      [8:0] n136;
wire      [8:0] n137;
wire            n138;
wire      [9:0] n139;
wire      [9:0] n140;
wire      [9:0] n141;
wire      [9:0] n142;
wire      [9:0] n143;
wire      [9:0] n144;
wire      [9:0] n145;
wire      [9:0] n146;
wire      [9:0] n147;
wire            n148;
wire    [647:0] n149;
wire      [7:0] n150;
wire      [7:0] n151;
wire      [7:0] n152;
wire      [7:0] n153;
wire      [7:0] n154;
wire      [7:0] n155;
wire      [7:0] n156;
wire            n157;
wire            n158;
wire            n159;
wire            n160;
wire            n161;
wire            n162;
wire            n163;
wire            n164;
wire            n165;
wire            n166;
wire            n167;
wire            n168;
wire            n169;
wire            n170;
wire     [18:0] n171;
wire            n172;
wire            n173;
wire            n174;
wire            n175;
wire            n176;
wire            n177;
wire            n178;
wire            n179;
wire            n180;
wire            n181;
wire            n182;
wire            n183;
wire            n184;
wire            n185;
wire            n186;
wire            n187;
wire            n188;
wire            n189;
wire            n190;
wire            n191;
wire            n192;
wire            n193;
wire            n194;
wire            n195;
wire            n196;
wire            n197;
wire            n198;
wire            n199;
wire            n200;
wire            n201;
wire            n202;
wire            n203;
wire            n204;
wire            n205;
wire            n206;
wire            n207;
wire            n208;
wire            n209;
wire            n210;
wire            n211;
wire            n212;
wire            n213;
wire            n214;
wire            n215;
wire            n216;
wire            n217;
wire            n218;
wire            n219;
wire            n220;
wire            n221;
wire            n222;
wire     [18:0] n223;
wire     [18:0] n224;
wire     [18:0] n225;
wire     [18:0] n226;
wire     [18:0] n227;
wire     [18:0] n228;
wire     [18:0] n229;
wire            n230;
wire            n231;
wire            n232;
wire            n233;
wire            n234;
wire            n235;
wire            n236;
wire            n237;
wire            n238;
wire            n239;
wire            n240;
wire            n241;
wire            n242;
wire            n243;
wire            n244;
wire            n245;
wire            n246;
wire            n247;
wire            n248;
wire            n249;
wire            n250;
wire            n251;
wire            n252;
wire            n253;
wire            n254;
wire            n255;
wire            n256;
wire            n257;
wire            n258;
wire            n259;
wire            n260;
wire            n261;
wire            n262;
wire            n263;
wire            n264;
wire            n265;
wire            n266;
wire            n267;
wire            n268;
wire            n269;
wire            n270;
wire            n271;
wire            n272;
wire            n273;
wire            n274;
wire            n275;
wire            n276;
wire            n277;
wire            n278;
wire            n279;
wire            n280;
wire            n281;
wire            n282;
wire            n283;
wire      [7:0] n284;
wire      [7:0] n285;
wire      [7:0] n286;
wire      [7:0] n287;
wire      [7:0] n288;
wire      [7:0] n289;
wire      [7:0] n290;
wire      [7:0] n291;
wire      [7:0] n292;
wire      [7:0] n293;
wire      [7:0] n294;
wire      [7:0] n295;
wire            n296;
wire            n297;
wire            n298;
wire            n299;
wire            n300;
wire            n301;
wire            n302;
wire            n303;
wire            n304;
wire            n305;
wire            n306;
wire            n307;
wire            n308;
wire            n309;
wire            n310;
wire            n311;
wire      [7:0] n312;
wire            n313;
wire      [7:0] n314;
wire            n315;
wire      [7:0] n316;
wire            n317;
wire      [7:0] n318;
wire            n319;
wire      [7:0] n320;
wire            n321;
wire      [7:0] n322;
wire            n323;
wire      [7:0] n324;
wire            n325;
wire      [7:0] n326;
wire      [7:0] n327;
wire      [7:0] n328;
wire      [7:0] n329;
wire      [7:0] n330;
wire      [7:0] n331;
wire      [7:0] n332;
wire      [7:0] n333;
wire      [7:0] n334;
wire      [7:0] n335;
wire      [7:0] n336;
wire      [7:0] n337;
wire      [7:0] n338;
wire      [7:0] n339;
wire      [7:0] n340;
wire      [7:0] n341;
wire      [7:0] n342;
wire      [7:0] n343;
wire      [7:0] n344;
wire      [7:0] n345;
wire      [7:0] n346;
wire      [7:0] n347;
wire      [7:0] n348;
wire      [7:0] n349;
wire      [7:0] n350;
wire      [7:0] n351;
wire      [7:0] n352;
wire      [7:0] n353;
wire      [7:0] n354;
wire      [7:0] n355;
wire      [7:0] n356;
wire      [7:0] n357;
wire      [7:0] n358;
wire      [7:0] n359;
wire      [7:0] n360;
wire      [7:0] n361;
wire      [7:0] n362;
wire      [7:0] n363;
wire      [7:0] n364;
wire      [7:0] n365;
wire      [7:0] n366;
wire      [7:0] n367;
wire      [7:0] n368;
wire      [7:0] n369;
wire      [7:0] n370;
wire      [7:0] n371;
wire      [7:0] n372;
wire      [7:0] n373;
wire      [7:0] n374;
wire      [7:0] n375;
wire      [7:0] n376;
wire      [7:0] n377;
wire      [7:0] n378;
wire      [7:0] n379;
wire      [7:0] n380;
wire      [7:0] n381;
wire      [7:0] n382;
wire      [7:0] n383;
wire     [15:0] n384;
wire     [23:0] n385;
wire     [31:0] n386;
wire     [39:0] n387;
wire     [47:0] n388;
wire     [55:0] n389;
wire     [63:0] n390;
wire     [71:0] n391;
wire     [71:0] n392;
wire     [71:0] n393;
wire     [71:0] n394;
wire     [71:0] n395;
wire     [71:0] n396;
wire     [71:0] n397;
wire     [71:0] n398;
wire     [71:0] n399;
wire     [71:0] n400;
wire     [71:0] n401;
wire     [71:0] n402;
wire     [71:0] n403;
wire     [71:0] n404;
wire     [71:0] n405;
wire            n406;
wire            n407;
wire            n408;
wire            n409;
wire            n410;
wire            n411;
wire            n412;
wire            n413;
wire            n414;
wire            n415;
wire            n416;
wire            n417;
wire            n418;
wire            n419;
wire            n420;
wire            n421;
wire            n422;
wire            n423;
wire      [7:0] n424;
wire      [7:0] n425;
wire      [7:0] n426;
wire      [7:0] n427;
wire      [7:0] n428;
wire      [7:0] n429;
wire      [7:0] n430;
wire      [7:0] n431;
wire      [7:0] n432;
wire     [15:0] n433;
wire     [23:0] n434;
wire     [31:0] n435;
wire     [39:0] n436;
wire     [47:0] n437;
wire     [55:0] n438;
wire     [63:0] n439;
wire     [71:0] n440;
wire      [7:0] n441;
wire      [7:0] n442;
wire      [7:0] n443;
wire      [7:0] n444;
wire      [7:0] n445;
wire      [7:0] n446;
wire      [7:0] n447;
wire      [7:0] n448;
wire      [7:0] n449;
wire     [15:0] n450;
wire     [23:0] n451;
wire     [31:0] n452;
wire     [39:0] n453;
wire     [47:0] n454;
wire     [55:0] n455;
wire     [63:0] n456;
wire     [71:0] n457;
wire      [7:0] n458;
wire      [7:0] n459;
wire      [7:0] n460;
wire      [7:0] n461;
wire      [7:0] n462;
wire      [7:0] n463;
wire      [7:0] n464;
wire      [7:0] n465;
wire      [7:0] n466;
wire     [15:0] n467;
wire     [23:0] n468;
wire     [31:0] n469;
wire     [39:0] n470;
wire     [47:0] n471;
wire     [55:0] n472;
wire     [63:0] n473;
wire     [71:0] n474;
wire      [7:0] n475;
wire      [7:0] n476;
wire      [7:0] n477;
wire      [7:0] n478;
wire      [7:0] n479;
wire      [7:0] n480;
wire      [7:0] n481;
wire      [7:0] n482;
wire      [7:0] n483;
wire     [15:0] n484;
wire     [23:0] n485;
wire     [31:0] n486;
wire     [39:0] n487;
wire     [47:0] n488;
wire     [55:0] n489;
wire     [63:0] n490;
wire     [71:0] n491;
wire      [7:0] n492;
wire      [7:0] n493;
wire      [7:0] n494;
wire      [7:0] n495;
wire      [7:0] n496;
wire      [7:0] n497;
wire      [7:0] n498;
wire      [7:0] n499;
wire      [7:0] n500;
wire     [15:0] n501;
wire     [23:0] n502;
wire     [31:0] n503;
wire     [39:0] n504;
wire     [47:0] n505;
wire     [55:0] n506;
wire     [63:0] n507;
wire     [71:0] n508;
wire      [7:0] n509;
wire      [7:0] n510;
wire      [7:0] n511;
wire      [7:0] n512;
wire      [7:0] n513;
wire      [7:0] n514;
wire      [7:0] n515;
wire      [7:0] n516;
wire      [7:0] n517;
wire     [15:0] n518;
wire     [23:0] n519;
wire     [31:0] n520;
wire     [39:0] n521;
wire     [47:0] n522;
wire     [55:0] n523;
wire     [63:0] n524;
wire     [71:0] n525;
wire      [7:0] n526;
wire      [7:0] n527;
wire      [7:0] n528;
wire      [7:0] n529;
wire      [7:0] n530;
wire      [7:0] n531;
wire      [7:0] n532;
wire      [7:0] n533;
wire      [7:0] n534;
wire     [15:0] n535;
wire     [23:0] n536;
wire     [31:0] n537;
wire     [39:0] n538;
wire     [47:0] n539;
wire     [55:0] n540;
wire     [63:0] n541;
wire     [71:0] n542;
wire      [7:0] n543;
wire      [7:0] n544;
wire      [7:0] n545;
wire      [7:0] n546;
wire      [7:0] n547;
wire      [7:0] n548;
wire      [7:0] n549;
wire      [7:0] n550;
wire      [7:0] n551;
wire     [15:0] n552;
wire     [23:0] n553;
wire     [31:0] n554;
wire     [39:0] n555;
wire     [47:0] n556;
wire     [55:0] n557;
wire     [63:0] n558;
wire     [71:0] n559;
wire      [7:0] n560;
wire      [7:0] n561;
wire      [7:0] n562;
wire      [7:0] n563;
wire      [7:0] n564;
wire      [7:0] n565;
wire      [7:0] n566;
wire      [7:0] n567;
wire      [7:0] n568;
wire     [15:0] n569;
wire     [23:0] n570;
wire     [31:0] n571;
wire     [39:0] n572;
wire     [47:0] n573;
wire     [55:0] n574;
wire     [63:0] n575;
wire     [71:0] n576;
wire    [143:0] n577;
wire    [215:0] n578;
wire    [287:0] n579;
wire    [359:0] n580;
wire    [431:0] n581;
wire    [503:0] n582;
wire    [575:0] n583;
wire    [647:0] n584;
wire    [647:0] n585;
wire    [647:0] n586;
wire    [647:0] n587;
wire    [647:0] n588;
wire    [647:0] n589;
wire    [647:0] n590;
wire    [647:0] n591;
wire    [647:0] n592;
wire    [647:0] n593;
wire    [647:0] n594;
wire    [647:0] n595;
wire    [647:0] n596;
wire    [647:0] n597;
wire            n598;
wire            n599;
wire            n600;
wire            n601;
wire            n602;
wire            n603;
wire            n604;
wire            n605;
wire            n606;
wire            n607;
wire            n608;
wire            n609;
wire            n610;
wire            n611;
wire            n612;
wire            n613;
wire            n614;
wire            n615;
wire      [8:0] LB2D_proc_0_addr0;
wire      [7:0] LB2D_proc_0_data0;
wire            n616;
wire            n617;
wire            n618;
wire            n619;
wire            n620;
wire            n621;
wire            n622;
wire            n623;
wire            n624;
wire            n625;
wire            n626;
wire            n627;
wire            n628;
wire            n629;
wire            n630;
wire            n631;
wire            n632;
wire            n633;
wire            n634;
wire      [8:0] LB2D_proc_1_addr0;
wire      [7:0] LB2D_proc_1_data0;
wire            n635;
wire            n636;
wire            n637;
wire      [8:0] LB2D_proc_2_addr0;
wire      [7:0] LB2D_proc_2_data0;
wire            n638;
wire            n639;
wire            n640;
wire      [8:0] LB2D_proc_3_addr0;
wire      [7:0] LB2D_proc_3_data0;
wire            n641;
wire            n642;
wire            n643;
wire      [8:0] LB2D_proc_4_addr0;
wire      [7:0] LB2D_proc_4_data0;
wire            n644;
wire            n645;
wire            n646;
wire      [8:0] LB2D_proc_5_addr0;
wire      [7:0] LB2D_proc_5_data0;
wire            n647;
wire            n648;
wire            n649;
wire      [8:0] LB2D_proc_6_addr0;
wire      [7:0] LB2D_proc_6_data0;
wire            n650;
wire            n651;
wire            n652;
wire      [8:0] LB2D_proc_7_addr0;
wire      [7:0] LB2D_proc_7_data0;
wire            n653;
wire            n654;
wire            n655;
wire            n656;
reg      [7:0] LB2D_proc_0[511:0];
reg      [7:0] LB2D_proc_1[511:0];
reg      [7:0] LB2D_proc_2[511:0];
reg      [7:0] LB2D_proc_3[511:0];
reg      [7:0] LB2D_proc_4[511:0];
reg      [7:0] LB2D_proc_5[511:0];
reg      [7:0] LB2D_proc_6[511:0];
reg      [7:0] LB2D_proc_7[511:0];
wire clk;
wire rst;
wire step;
assign n0 =  ( arg_0_TREADY ) == ( 1'd1 )  ;
assign n1 =  ( arg_0_TVALID ) == ( 1'd1 )  ;
assign n2 =  ( n0 ) & ( n1 )  ;
assign n3 =  ( arg_1_TVALID ) == ( 1'd0 )  ;
assign n4 =  ( n2 ) & ( n3 )  ;
assign n5 =  ( arg_1_TREADY ) == ( 1'd1 )  ;
assign n6 =  ( arg_1_TVALID ) == ( 1'd1 )  ;
assign n7 =  ( n5 ) & ( n6 )  ;
assign n8 =  ( arg_0_TREADY ) == ( 1'd0 )  ;
assign n9 =  ( n7 ) & ( n8 )  ;
assign n10 =  ( arg_0_TVALID ) == ( 1'd0 )  ;
assign n11 =  ( gb_exit_it_1 ) == ( 1'd0 )  ;
assign n12 =  ( stencil_stream_empty ) == ( 1'd0 )  ;
assign n13 =  ( n11 ) & ( n12 )  ;
assign n14 =  ( gb_exit_it_1 ) == ( 1'd1 )  ;
assign n15 =  ( gb_exit_it_8 ) == ( 1'd0 )  ;
assign n16 =  ( n14 ) & ( n15 )  ;
assign n17 =  ( n13 ) | ( n16 )  ;
assign n18 =  ( n10 ) & ( n17 )  ;
assign n19 =  ( slice_stream_empty ) == ( 1'd0 )  ;
assign n20 =  ( stencil_stream_full ) == ( 1'd0 )  ;
assign n21 =  ( LB2D_shift_x ) < ( 9'd8 )  ;
assign n22 =  ( n20 ) | ( n21 )  ;
assign n23 =  ( n19 ) & ( n22 )  ;
assign n24 =  ( in_stream_empty ) == ( 1'd0 )  ;
assign n25 =  ( LB2D_proc_x ) != ( 9'd488 )  ;
assign n26 =  ( n24 ) & ( n25 )  ;
assign n27 =  ( slice_stream_full ) == ( 1'd0 )  ;
assign n28 =  ( LB2D_proc_y ) < ( 10'd8 )  ;
assign n29 =  ( n27 ) | ( n28 )  ;
assign n30 =  ( n26 ) & ( n29 )  ;
assign n31 =  ( arg_1_TREADY ) == ( 1'd0 )  ;
assign n32 =  ( in_stream_full ) == ( 1'd0 )  ;
assign n33 =  ( n31 ) & ( n32 )  ;
assign n34 =  ( LB1D_p_cnt ) != ( 19'd316224 )  ;
assign n35 =  ( n33 ) & ( n34 )  ;
assign n36 =  ( n35 ) ? ( LB1D_buff ) : ( LB1D_buff ) ;
assign n37 =  ( n30 ) ? ( LB1D_buff ) : ( n36 ) ;
assign n38 =  ( n23 ) ? ( LB1D_buff ) : ( n37 ) ;
assign n39 =  ( n18 ) ? ( LB1D_buff ) : ( n38 ) ;
assign n40 =  ( n9 ) ? ( arg_1_TDATA ) : ( n39 ) ;
assign n41 =  ( n4 ) ? ( arg_1_TDATA ) : ( n40 ) ;
assign n42 =  ( LB1D_p_cnt ) + ( 19'd1 )  ;
assign n43 =  ( n35 ) ? ( n42 ) : ( LB1D_p_cnt ) ;
assign n44 =  ( n30 ) ? ( LB1D_p_cnt ) : ( n43 ) ;
assign n45 =  ( n23 ) ? ( LB1D_p_cnt ) : ( n44 ) ;
assign n46 =  ( n18 ) ? ( LB1D_p_cnt ) : ( n45 ) ;
assign n47 =  ( n9 ) ? ( LB1D_p_cnt ) : ( n46 ) ;
assign n48 =  ( n4 ) ? ( LB1D_p_cnt ) : ( n47 ) ;
assign n49 =  ( LB2D_proc_w ) < ( 64'd7 )  ;
assign n50 =  ( LB2D_proc_x ) < ( 9'd488 )  ;
assign n51 =  ( LB2D_proc_w ) + ( 64'd1 )  ;
assign n52 =  ( n50 ) ? ( LB2D_proc_w ) : ( n51 ) ;
assign n53 =  ( n49 ) ? ( n52 ) : ( 64'd0 ) ;
assign n54 =  ( n35 ) ? ( LB2D_proc_w ) : ( LB2D_proc_w ) ;
assign n55 =  ( n30 ) ? ( n53 ) : ( n54 ) ;
assign n56 =  ( n23 ) ? ( LB2D_proc_w ) : ( n55 ) ;
assign n57 =  ( n18 ) ? ( LB2D_proc_w ) : ( n56 ) ;
assign n58 =  ( n9 ) ? ( LB2D_proc_w ) : ( n57 ) ;
assign n59 =  ( n4 ) ? ( LB2D_proc_w ) : ( n58 ) ;
assign n60 =  ( LB2D_proc_x ) == ( 9'd488 )  ;
assign n61 =  ( n24 ) & ( n60 )  ;
assign n62 =  ( n61 ) & ( n29 )  ;
assign n63 =  ( LB2D_proc_x ) + ( 9'd1 )  ;
assign n64 =  ( n35 ) ? ( LB2D_proc_x ) : ( LB2D_proc_x ) ;
assign n65 =  ( n30 ) ? ( n63 ) : ( n64 ) ;
assign n66 =  ( n62 ) ? ( 9'd0 ) : ( n65 ) ;
assign n67 =  ( n23 ) ? ( LB2D_proc_x ) : ( n66 ) ;
assign n68 =  ( n18 ) ? ( LB2D_proc_x ) : ( n67 ) ;
assign n69 =  ( n9 ) ? ( LB2D_proc_x ) : ( n68 ) ;
assign n70 =  ( n4 ) ? ( LB2D_proc_x ) : ( n69 ) ;
assign n71 =  ( LB2D_proc_y ) < ( 10'd488 )  ;
assign n72 =  ( n71 ) ? ( LB2D_proc_y ) : ( 10'd488 ) ;
assign n73 =  ( n35 ) ? ( LB2D_proc_y ) : ( LB2D_proc_y ) ;
assign n74 =  ( n30 ) ? ( n72 ) : ( n73 ) ;
assign n75 =  ( n23 ) ? ( LB2D_proc_y ) : ( n74 ) ;
assign n76 =  ( n18 ) ? ( LB2D_proc_y ) : ( n75 ) ;
assign n77 =  ( n9 ) ? ( LB2D_proc_y ) : ( n76 ) ;
assign n78 =  ( n4 ) ? ( LB2D_proc_y ) : ( n77 ) ;
assign n79 =  ( slice_stream_full ) == ( 1'd1 )  ;
assign n80 =  ( n79 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n81 =  ( n35 ) ? ( LB2D_shift_0 ) : ( LB2D_shift_0 ) ;
assign n82 =  ( n30 ) ? ( LB2D_shift_0 ) : ( n81 ) ;
assign n83 =  ( n23 ) ? ( n80 ) : ( n82 ) ;
assign n84 =  ( n18 ) ? ( LB2D_shift_0 ) : ( n83 ) ;
assign n85 =  ( n9 ) ? ( LB2D_shift_0 ) : ( n84 ) ;
assign n86 =  ( n4 ) ? ( LB2D_shift_0 ) : ( n85 ) ;
assign n87 =  ( n35 ) ? ( LB2D_shift_1 ) : ( LB2D_shift_1 ) ;
assign n88 =  ( n30 ) ? ( LB2D_shift_1 ) : ( n87 ) ;
assign n89 =  ( n23 ) ? ( LB2D_shift_0 ) : ( n88 ) ;
assign n90 =  ( n18 ) ? ( LB2D_shift_1 ) : ( n89 ) ;
assign n91 =  ( n9 ) ? ( LB2D_shift_1 ) : ( n90 ) ;
assign n92 =  ( n4 ) ? ( LB2D_shift_1 ) : ( n91 ) ;
assign n93 =  ( n35 ) ? ( LB2D_shift_2 ) : ( LB2D_shift_2 ) ;
assign n94 =  ( n30 ) ? ( LB2D_shift_2 ) : ( n93 ) ;
assign n95 =  ( n23 ) ? ( LB2D_shift_1 ) : ( n94 ) ;
assign n96 =  ( n18 ) ? ( LB2D_shift_2 ) : ( n95 ) ;
assign n97 =  ( n9 ) ? ( LB2D_shift_2 ) : ( n96 ) ;
assign n98 =  ( n4 ) ? ( LB2D_shift_2 ) : ( n97 ) ;
assign n99 =  ( n35 ) ? ( LB2D_shift_3 ) : ( LB2D_shift_3 ) ;
assign n100 =  ( n30 ) ? ( LB2D_shift_3 ) : ( n99 ) ;
assign n101 =  ( n23 ) ? ( LB2D_shift_2 ) : ( n100 ) ;
assign n102 =  ( n18 ) ? ( LB2D_shift_3 ) : ( n101 ) ;
assign n103 =  ( n9 ) ? ( LB2D_shift_3 ) : ( n102 ) ;
assign n104 =  ( n4 ) ? ( LB2D_shift_3 ) : ( n103 ) ;
assign n105 =  ( n35 ) ? ( LB2D_shift_4 ) : ( LB2D_shift_4 ) ;
assign n106 =  ( n30 ) ? ( LB2D_shift_4 ) : ( n105 ) ;
assign n107 =  ( n23 ) ? ( LB2D_shift_3 ) : ( n106 ) ;
assign n108 =  ( n18 ) ? ( LB2D_shift_4 ) : ( n107 ) ;
assign n109 =  ( n9 ) ? ( LB2D_shift_4 ) : ( n108 ) ;
assign n110 =  ( n4 ) ? ( LB2D_shift_4 ) : ( n109 ) ;
assign n111 =  ( n35 ) ? ( LB2D_shift_5 ) : ( LB2D_shift_5 ) ;
assign n112 =  ( n30 ) ? ( LB2D_shift_5 ) : ( n111 ) ;
assign n113 =  ( n23 ) ? ( LB2D_shift_4 ) : ( n112 ) ;
assign n114 =  ( n18 ) ? ( LB2D_shift_5 ) : ( n113 ) ;
assign n115 =  ( n9 ) ? ( LB2D_shift_5 ) : ( n114 ) ;
assign n116 =  ( n4 ) ? ( LB2D_shift_5 ) : ( n115 ) ;
assign n117 =  ( n35 ) ? ( LB2D_shift_6 ) : ( LB2D_shift_6 ) ;
assign n118 =  ( n30 ) ? ( LB2D_shift_6 ) : ( n117 ) ;
assign n119 =  ( n23 ) ? ( LB2D_shift_5 ) : ( n118 ) ;
assign n120 =  ( n18 ) ? ( LB2D_shift_6 ) : ( n119 ) ;
assign n121 =  ( n9 ) ? ( LB2D_shift_6 ) : ( n120 ) ;
assign n122 =  ( n4 ) ? ( LB2D_shift_6 ) : ( n121 ) ;
assign n123 =  ( n35 ) ? ( LB2D_shift_7 ) : ( LB2D_shift_7 ) ;
assign n124 =  ( n30 ) ? ( LB2D_shift_7 ) : ( n123 ) ;
assign n125 =  ( n23 ) ? ( LB2D_shift_6 ) : ( n124 ) ;
assign n126 =  ( n18 ) ? ( LB2D_shift_7 ) : ( n125 ) ;
assign n127 =  ( n9 ) ? ( LB2D_shift_7 ) : ( n126 ) ;
assign n128 =  ( n4 ) ? ( LB2D_shift_7 ) : ( n127 ) ;
assign n129 =  ( LB2D_shift_x ) < ( 9'd487 )  ;
assign n130 =  ( LB2D_shift_x ) + ( 9'd1 )  ;
assign n131 =  ( n129 ) ? ( n130 ) : ( 9'd0 ) ;
assign n132 =  ( n35 ) ? ( LB2D_shift_x ) : ( LB2D_shift_x ) ;
assign n133 =  ( n30 ) ? ( LB2D_shift_x ) : ( n132 ) ;
assign n134 =  ( n23 ) ? ( n131 ) : ( n133 ) ;
assign n135 =  ( n18 ) ? ( LB2D_shift_x ) : ( n134 ) ;
assign n136 =  ( n9 ) ? ( LB2D_shift_x ) : ( n135 ) ;
assign n137 =  ( n4 ) ? ( LB2D_shift_x ) : ( n136 ) ;
assign n138 =  ( LB2D_shift_y ) < ( 10'd479 )  ;
assign n139 =  ( LB2D_shift_y ) + ( 10'd1 )  ;
assign n140 =  ( n129 ) ? ( LB2D_shift_y ) : ( n139 ) ;
assign n141 =  ( n138 ) ? ( n140 ) : ( 10'd479 ) ;
assign n142 =  ( n35 ) ? ( LB2D_shift_y ) : ( LB2D_shift_y ) ;
assign n143 =  ( n30 ) ? ( LB2D_shift_y ) : ( n142 ) ;
assign n144 =  ( n23 ) ? ( n141 ) : ( n143 ) ;
assign n145 =  ( n18 ) ? ( LB2D_shift_y ) : ( n144 ) ;
assign n146 =  ( n9 ) ? ( LB2D_shift_y ) : ( n145 ) ;
assign n147 =  ( n4 ) ? ( LB2D_shift_y ) : ( n146 ) ;
assign n148 =  ( stencil_stream_full ) == ( 1'd1 )  ;
assign n149 =  ( n148 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_0 ) ;
//assign n150 = gb_fun(n149) ;
gb_fun gb_fun_U (
    .stencil (n149),
    .result (n150)
);

assign n151 =  ( n35 ) ? ( arg_0_TDATA ) : ( arg_0_TDATA ) ;
assign n152 =  ( n30 ) ? ( arg_0_TDATA ) : ( n151 ) ;
assign n153 =  ( n23 ) ? ( arg_0_TDATA ) : ( n152 ) ;
assign n154 =  ( n18 ) ? ( n150 ) : ( n153 ) ;
assign n155 =  ( n9 ) ? ( arg_0_TDATA ) : ( n154 ) ;
assign n156 =  ( n4 ) ? ( arg_0_TDATA ) : ( n155 ) ;
assign n157 =  ( gb_pp_it_8 ) == ( 1'd1 )  ;
assign n158 =  ( n157 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n159 =  ( n35 ) ? ( arg_0_TVALID ) : ( arg_0_TVALID ) ;
assign n160 =  ( n30 ) ? ( arg_0_TVALID ) : ( n159 ) ;
assign n161 =  ( n23 ) ? ( arg_0_TVALID ) : ( n160 ) ;
assign n162 =  ( n18 ) ? ( n158 ) : ( n161 ) ;
assign n163 =  ( n9 ) ? ( arg_0_TVALID ) : ( n162 ) ;
assign n164 =  ( n4 ) ? ( 1'd0 ) : ( n163 ) ;
assign n165 =  ( n35 ) ? ( 1'd1 ) : ( arg_1_TREADY ) ;
assign n166 =  ( n30 ) ? ( arg_1_TREADY ) : ( n165 ) ;
assign n167 =  ( n23 ) ? ( arg_1_TREADY ) : ( n166 ) ;
assign n168 =  ( n18 ) ? ( arg_1_TREADY ) : ( n167 ) ;
assign n169 =  ( n9 ) ? ( 1'd0 ) : ( n168 ) ;
assign n170 =  ( n4 ) ? ( 1'd0 ) : ( n169 ) ;
assign n171 =  ( gb_p_cnt ) + ( 19'd1 )  ;
assign n172 =  ( n171 ) == ( 19'd307200 )  ;
assign n173 =  ( n172 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n174 =  ( n35 ) ? ( gb_exit_it_1 ) : ( gb_exit_it_1 ) ;
assign n175 =  ( n30 ) ? ( gb_exit_it_1 ) : ( n174 ) ;
assign n176 =  ( n23 ) ? ( gb_exit_it_1 ) : ( n175 ) ;
assign n177 =  ( n18 ) ? ( n173 ) : ( n176 ) ;
assign n178 =  ( n9 ) ? ( gb_exit_it_1 ) : ( n177 ) ;
assign n179 =  ( n4 ) ? ( gb_exit_it_1 ) : ( n178 ) ;
assign n180 =  ( n35 ) ? ( gb_exit_it_2 ) : ( gb_exit_it_2 ) ;
assign n181 =  ( n30 ) ? ( gb_exit_it_2 ) : ( n180 ) ;
assign n182 =  ( n23 ) ? ( gb_exit_it_2 ) : ( n181 ) ;
assign n183 =  ( n18 ) ? ( gb_exit_it_1 ) : ( n182 ) ;
assign n184 =  ( n9 ) ? ( gb_exit_it_2 ) : ( n183 ) ;
assign n185 =  ( n4 ) ? ( gb_exit_it_2 ) : ( n184 ) ;
assign n186 =  ( n35 ) ? ( gb_exit_it_3 ) : ( gb_exit_it_3 ) ;
assign n187 =  ( n30 ) ? ( gb_exit_it_3 ) : ( n186 ) ;
assign n188 =  ( n23 ) ? ( gb_exit_it_3 ) : ( n187 ) ;
assign n189 =  ( n18 ) ? ( gb_exit_it_2 ) : ( n188 ) ;
assign n190 =  ( n9 ) ? ( gb_exit_it_3 ) : ( n189 ) ;
assign n191 =  ( n4 ) ? ( gb_exit_it_3 ) : ( n190 ) ;
assign n192 =  ( n35 ) ? ( gb_exit_it_4 ) : ( gb_exit_it_4 ) ;
assign n193 =  ( n30 ) ? ( gb_exit_it_4 ) : ( n192 ) ;
assign n194 =  ( n23 ) ? ( gb_exit_it_4 ) : ( n193 ) ;
assign n195 =  ( n18 ) ? ( gb_exit_it_3 ) : ( n194 ) ;
assign n196 =  ( n9 ) ? ( gb_exit_it_4 ) : ( n195 ) ;
assign n197 =  ( n4 ) ? ( gb_exit_it_4 ) : ( n196 ) ;
assign n198 =  ( n35 ) ? ( gb_exit_it_5 ) : ( gb_exit_it_5 ) ;
assign n199 =  ( n30 ) ? ( gb_exit_it_5 ) : ( n198 ) ;
assign n200 =  ( n23 ) ? ( gb_exit_it_5 ) : ( n199 ) ;
assign n201 =  ( n18 ) ? ( gb_exit_it_4 ) : ( n200 ) ;
assign n202 =  ( n9 ) ? ( gb_exit_it_5 ) : ( n201 ) ;
assign n203 =  ( n4 ) ? ( gb_exit_it_5 ) : ( n202 ) ;
assign n204 =  ( n35 ) ? ( gb_exit_it_6 ) : ( gb_exit_it_6 ) ;
assign n205 =  ( n30 ) ? ( gb_exit_it_6 ) : ( n204 ) ;
assign n206 =  ( n23 ) ? ( gb_exit_it_6 ) : ( n205 ) ;
assign n207 =  ( n18 ) ? ( gb_exit_it_5 ) : ( n206 ) ;
assign n208 =  ( n9 ) ? ( gb_exit_it_6 ) : ( n207 ) ;
assign n209 =  ( n4 ) ? ( gb_exit_it_6 ) : ( n208 ) ;
assign n210 =  ( n35 ) ? ( gb_exit_it_7 ) : ( gb_exit_it_7 ) ;
assign n211 =  ( n30 ) ? ( gb_exit_it_7 ) : ( n210 ) ;
assign n212 =  ( n23 ) ? ( gb_exit_it_7 ) : ( n211 ) ;
assign n213 =  ( n18 ) ? ( gb_exit_it_6 ) : ( n212 ) ;
assign n214 =  ( n9 ) ? ( gb_exit_it_7 ) : ( n213 ) ;
assign n215 =  ( n4 ) ? ( gb_exit_it_7 ) : ( n214 ) ;
assign n216 =  ( n35 ) ? ( gb_exit_it_8 ) : ( gb_exit_it_8 ) ;
assign n217 =  ( n30 ) ? ( gb_exit_it_8 ) : ( n216 ) ;
assign n218 =  ( n23 ) ? ( gb_exit_it_8 ) : ( n217 ) ;
assign n219 =  ( n18 ) ? ( gb_exit_it_7 ) : ( n218 ) ;
assign n220 =  ( n9 ) ? ( gb_exit_it_8 ) : ( n219 ) ;
assign n221 =  ( n4 ) ? ( gb_exit_it_8 ) : ( n220 ) ;
assign n222 =  ( gb_p_cnt ) < ( 19'd307200 )  ;
assign n223 =  ( n222 ) ? ( n171 ) : ( 19'd307200 ) ;
assign n224 =  ( n35 ) ? ( gb_p_cnt ) : ( gb_p_cnt ) ;
assign n225 =  ( n30 ) ? ( gb_p_cnt ) : ( n224 ) ;
assign n226 =  ( n23 ) ? ( gb_p_cnt ) : ( n225 ) ;
assign n227 =  ( n18 ) ? ( n223 ) : ( n226 ) ;
assign n228 =  ( n9 ) ? ( gb_p_cnt ) : ( n227 ) ;
assign n229 =  ( n4 ) ? ( gb_p_cnt ) : ( n228 ) ;
assign n230 =  ( n35 ) ? ( gb_pp_it_1 ) : ( gb_pp_it_1 ) ;
assign n231 =  ( n30 ) ? ( gb_pp_it_1 ) : ( n230 ) ;
assign n232 =  ( n23 ) ? ( gb_pp_it_1 ) : ( n231 ) ;
assign n233 =  ( n18 ) ? ( 1'd1 ) : ( n232 ) ;
assign n234 =  ( n9 ) ? ( gb_pp_it_1 ) : ( n233 ) ;
assign n235 =  ( n4 ) ? ( gb_pp_it_1 ) : ( n234 ) ;
assign n236 =  ( n35 ) ? ( gb_pp_it_2 ) : ( gb_pp_it_2 ) ;
assign n237 =  ( n30 ) ? ( gb_pp_it_2 ) : ( n236 ) ;
assign n238 =  ( n23 ) ? ( gb_pp_it_2 ) : ( n237 ) ;
assign n239 =  ( n18 ) ? ( gb_pp_it_1 ) : ( n238 ) ;
assign n240 =  ( n9 ) ? ( gb_pp_it_2 ) : ( n239 ) ;
assign n241 =  ( n4 ) ? ( gb_pp_it_2 ) : ( n240 ) ;
assign n242 =  ( n35 ) ? ( gb_pp_it_3 ) : ( gb_pp_it_3 ) ;
assign n243 =  ( n30 ) ? ( gb_pp_it_3 ) : ( n242 ) ;
assign n244 =  ( n23 ) ? ( gb_pp_it_3 ) : ( n243 ) ;
assign n245 =  ( n18 ) ? ( gb_pp_it_2 ) : ( n244 ) ;
assign n246 =  ( n9 ) ? ( gb_pp_it_3 ) : ( n245 ) ;
assign n247 =  ( n4 ) ? ( gb_pp_it_3 ) : ( n246 ) ;
assign n248 =  ( n35 ) ? ( gb_pp_it_4 ) : ( gb_pp_it_4 ) ;
assign n249 =  ( n30 ) ? ( gb_pp_it_4 ) : ( n248 ) ;
assign n250 =  ( n23 ) ? ( gb_pp_it_4 ) : ( n249 ) ;
assign n251 =  ( n18 ) ? ( gb_pp_it_3 ) : ( n250 ) ;
assign n252 =  ( n9 ) ? ( gb_pp_it_4 ) : ( n251 ) ;
assign n253 =  ( n4 ) ? ( gb_pp_it_4 ) : ( n252 ) ;
assign n254 =  ( n35 ) ? ( gb_pp_it_5 ) : ( gb_pp_it_5 ) ;
assign n255 =  ( n30 ) ? ( gb_pp_it_5 ) : ( n254 ) ;
assign n256 =  ( n23 ) ? ( gb_pp_it_5 ) : ( n255 ) ;
assign n257 =  ( n18 ) ? ( gb_pp_it_4 ) : ( n256 ) ;
assign n258 =  ( n9 ) ? ( gb_pp_it_5 ) : ( n257 ) ;
assign n259 =  ( n4 ) ? ( gb_pp_it_5 ) : ( n258 ) ;
assign n260 =  ( n35 ) ? ( gb_pp_it_6 ) : ( gb_pp_it_6 ) ;
assign n261 =  ( n30 ) ? ( gb_pp_it_6 ) : ( n260 ) ;
assign n262 =  ( n23 ) ? ( gb_pp_it_6 ) : ( n261 ) ;
assign n263 =  ( n18 ) ? ( gb_pp_it_5 ) : ( n262 ) ;
assign n264 =  ( n9 ) ? ( gb_pp_it_6 ) : ( n263 ) ;
assign n265 =  ( n4 ) ? ( gb_pp_it_6 ) : ( n264 ) ;
assign n266 =  ( n35 ) ? ( gb_pp_it_7 ) : ( gb_pp_it_7 ) ;
assign n267 =  ( n30 ) ? ( gb_pp_it_7 ) : ( n266 ) ;
assign n268 =  ( n23 ) ? ( gb_pp_it_7 ) : ( n267 ) ;
assign n269 =  ( n18 ) ? ( gb_pp_it_6 ) : ( n268 ) ;
assign n270 =  ( n9 ) ? ( gb_pp_it_7 ) : ( n269 ) ;
assign n271 =  ( n4 ) ? ( gb_pp_it_7 ) : ( n270 ) ;
assign n272 =  ( n35 ) ? ( gb_pp_it_8 ) : ( gb_pp_it_8 ) ;
assign n273 =  ( n30 ) ? ( gb_pp_it_8 ) : ( n272 ) ;
assign n274 =  ( n23 ) ? ( gb_pp_it_8 ) : ( n273 ) ;
assign n275 =  ( n18 ) ? ( gb_pp_it_7 ) : ( n274 ) ;
assign n276 =  ( n9 ) ? ( gb_pp_it_8 ) : ( n275 ) ;
assign n277 =  ( n4 ) ? ( gb_pp_it_8 ) : ( n276 ) ;
assign n278 =  ( n35 ) ? ( gb_pp_it_9 ) : ( gb_pp_it_9 ) ;
assign n279 =  ( n30 ) ? ( gb_pp_it_9 ) : ( n278 ) ;
assign n280 =  ( n23 ) ? ( gb_pp_it_9 ) : ( n279 ) ;
assign n281 =  ( n18 ) ? ( gb_pp_it_8 ) : ( n280 ) ;
assign n282 =  ( n9 ) ? ( gb_pp_it_9 ) : ( n281 ) ;
assign n283 =  ( n4 ) ? ( gb_pp_it_9 ) : ( n282 ) ;
assign n284 =  ( n35 ) ? ( LB1D_buff ) : ( in_stream_buff_0 ) ;
assign n285 =  ( n30 ) ? ( in_stream_buff_0 ) : ( n284 ) ;
assign n286 =  ( n23 ) ? ( in_stream_buff_0 ) : ( n285 ) ;
assign n287 =  ( n18 ) ? ( in_stream_buff_0 ) : ( n286 ) ;
assign n288 =  ( n9 ) ? ( in_stream_buff_0 ) : ( n287 ) ;
assign n289 =  ( n4 ) ? ( in_stream_buff_0 ) : ( n288 ) ;
assign n290 =  ( n35 ) ? ( in_stream_buff_0 ) : ( in_stream_buff_1 ) ;
assign n291 =  ( n30 ) ? ( in_stream_buff_1 ) : ( n290 ) ;
assign n292 =  ( n23 ) ? ( in_stream_buff_1 ) : ( n291 ) ;
assign n293 =  ( n18 ) ? ( in_stream_buff_1 ) : ( n292 ) ;
assign n294 =  ( n9 ) ? ( in_stream_buff_1 ) : ( n293 ) ;
assign n295 =  ( n4 ) ? ( in_stream_buff_1 ) : ( n294 ) ;
assign n296 =  ( in_stream_full ) == ( 1'd1 )  ;
assign n297 =  ( n296 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n298 =  ( n35 ) ? ( 1'd0 ) : ( in_stream_empty ) ;
assign n299 =  ( n30 ) ? ( n297 ) : ( n298 ) ;
assign n300 =  ( n23 ) ? ( in_stream_empty ) : ( n299 ) ;
assign n301 =  ( n18 ) ? ( in_stream_empty ) : ( n300 ) ;
assign n302 =  ( n9 ) ? ( in_stream_empty ) : ( n301 ) ;
assign n303 =  ( n4 ) ? ( in_stream_empty ) : ( n302 ) ;
assign n304 =  ( in_stream_empty ) == ( 1'd1 )  ;
assign n305 =  ( n304 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n306 =  ( n35 ) ? ( n305 ) : ( in_stream_full ) ;
assign n307 =  ( n30 ) ? ( 1'd0 ) : ( n306 ) ;
assign n308 =  ( n23 ) ? ( in_stream_full ) : ( n307 ) ;
assign n309 =  ( n18 ) ? ( in_stream_full ) : ( n308 ) ;
assign n310 =  ( n9 ) ? ( in_stream_full ) : ( n309 ) ;
assign n311 =  ( n4 ) ? ( in_stream_full ) : ( n310 ) ;
assign n312 =  ( n296 ) ? ( in_stream_buff_1 ) : ( in_stream_buff_0 ) ;
assign n313 =  ( LB2D_proc_w ) == ( 64'd0 )  ;
assign n314 =  (  LB2D_proc_7 [ LB2D_proc_x ] )  ;
assign n315 =  ( LB2D_proc_w ) == ( 64'd1 )  ;
assign n316 =  (  LB2D_proc_0 [ LB2D_proc_x ] )  ;
assign n317 =  ( LB2D_proc_w ) == ( 64'd2 )  ;
assign n318 =  (  LB2D_proc_1 [ LB2D_proc_x ] )  ;
assign n319 =  ( LB2D_proc_w ) == ( 64'd3 )  ;
assign n320 =  (  LB2D_proc_2 [ LB2D_proc_x ] )  ;
assign n321 =  ( LB2D_proc_w ) == ( 64'd4 )  ;
assign n322 =  (  LB2D_proc_3 [ LB2D_proc_x ] )  ;
assign n323 =  ( LB2D_proc_w ) == ( 64'd5 )  ;
assign n324 =  (  LB2D_proc_4 [ LB2D_proc_x ] )  ;
assign n325 =  ( LB2D_proc_w ) == ( 64'd6 )  ;
assign n326 =  (  LB2D_proc_5 [ LB2D_proc_x ] )  ;
assign n327 =  (  LB2D_proc_6 [ LB2D_proc_x ] )  ;
assign n328 =  ( n325 ) ? ( n326 ) : ( n327 ) ;
assign n329 =  ( n323 ) ? ( n324 ) : ( n328 ) ;
assign n330 =  ( n321 ) ? ( n322 ) : ( n329 ) ;
assign n331 =  ( n319 ) ? ( n320 ) : ( n330 ) ;
assign n332 =  ( n317 ) ? ( n318 ) : ( n331 ) ;
assign n333 =  ( n315 ) ? ( n316 ) : ( n332 ) ;
assign n334 =  ( n313 ) ? ( n314 ) : ( n333 ) ;
assign n335 =  ( n325 ) ? ( n324 ) : ( n326 ) ;
assign n336 =  ( n323 ) ? ( n322 ) : ( n335 ) ;
assign n337 =  ( n321 ) ? ( n320 ) : ( n336 ) ;
assign n338 =  ( n319 ) ? ( n318 ) : ( n337 ) ;
assign n339 =  ( n317 ) ? ( n316 ) : ( n338 ) ;
assign n340 =  ( n315 ) ? ( n314 ) : ( n339 ) ;
assign n341 =  ( n313 ) ? ( n327 ) : ( n340 ) ;
assign n342 =  ( n325 ) ? ( n322 ) : ( n324 ) ;
assign n343 =  ( n323 ) ? ( n320 ) : ( n342 ) ;
assign n344 =  ( n321 ) ? ( n318 ) : ( n343 ) ;
assign n345 =  ( n319 ) ? ( n316 ) : ( n344 ) ;
assign n346 =  ( n317 ) ? ( n314 ) : ( n345 ) ;
assign n347 =  ( n315 ) ? ( n327 ) : ( n346 ) ;
assign n348 =  ( n313 ) ? ( n326 ) : ( n347 ) ;
assign n349 =  ( n325 ) ? ( n320 ) : ( n322 ) ;
assign n350 =  ( n323 ) ? ( n318 ) : ( n349 ) ;
assign n351 =  ( n321 ) ? ( n316 ) : ( n350 ) ;
assign n352 =  ( n319 ) ? ( n314 ) : ( n351 ) ;
assign n353 =  ( n317 ) ? ( n327 ) : ( n352 ) ;
assign n354 =  ( n315 ) ? ( n326 ) : ( n353 ) ;
assign n355 =  ( n313 ) ? ( n324 ) : ( n354 ) ;
assign n356 =  ( n325 ) ? ( n318 ) : ( n320 ) ;
assign n357 =  ( n323 ) ? ( n316 ) : ( n356 ) ;
assign n358 =  ( n321 ) ? ( n314 ) : ( n357 ) ;
assign n359 =  ( n319 ) ? ( n327 ) : ( n358 ) ;
assign n360 =  ( n317 ) ? ( n326 ) : ( n359 ) ;
assign n361 =  ( n315 ) ? ( n324 ) : ( n360 ) ;
assign n362 =  ( n313 ) ? ( n322 ) : ( n361 ) ;
assign n363 =  ( n325 ) ? ( n316 ) : ( n318 ) ;
assign n364 =  ( n323 ) ? ( n314 ) : ( n363 ) ;
assign n365 =  ( n321 ) ? ( n327 ) : ( n364 ) ;
assign n366 =  ( n319 ) ? ( n326 ) : ( n365 ) ;
assign n367 =  ( n317 ) ? ( n324 ) : ( n366 ) ;
assign n368 =  ( n315 ) ? ( n322 ) : ( n367 ) ;
assign n369 =  ( n313 ) ? ( n320 ) : ( n368 ) ;
assign n370 =  ( n325 ) ? ( n314 ) : ( n316 ) ;
assign n371 =  ( n323 ) ? ( n327 ) : ( n370 ) ;
assign n372 =  ( n321 ) ? ( n326 ) : ( n371 ) ;
assign n373 =  ( n319 ) ? ( n324 ) : ( n372 ) ;
assign n374 =  ( n317 ) ? ( n322 ) : ( n373 ) ;
assign n375 =  ( n315 ) ? ( n320 ) : ( n374 ) ;
assign n376 =  ( n313 ) ? ( n318 ) : ( n375 ) ;
assign n377 =  ( n325 ) ? ( n327 ) : ( n314 ) ;
assign n378 =  ( n323 ) ? ( n326 ) : ( n377 ) ;
assign n379 =  ( n321 ) ? ( n324 ) : ( n378 ) ;
assign n380 =  ( n319 ) ? ( n322 ) : ( n379 ) ;
assign n381 =  ( n317 ) ? ( n320 ) : ( n380 ) ;
assign n382 =  ( n315 ) ? ( n318 ) : ( n381 ) ;
assign n383 =  ( n313 ) ? ( n316 ) : ( n382 ) ;
assign n384 =  { ( n376 ) , ( n383 ) }  ;
assign n385 =  { ( n369 ) , ( n384 ) }  ;
assign n386 =  { ( n362 ) , ( n385 ) }  ;
assign n387 =  { ( n355 ) , ( n386 ) }  ;
assign n388 =  { ( n348 ) , ( n387 ) }  ;
assign n389 =  { ( n341 ) , ( n388 ) }  ;
assign n390 =  { ( n334 ) , ( n389 ) }  ;
assign n391 =  { ( n312 ) , ( n390 ) }  ;
assign n392 =  ( n28 ) ? ( slice_stream_buff_0 ) : ( n391 ) ;
assign n393 =  ( n35 ) ? ( slice_stream_buff_0 ) : ( slice_stream_buff_0 ) ;
assign n394 =  ( n30 ) ? ( n392 ) : ( n393 ) ;
assign n395 =  ( n23 ) ? ( slice_stream_buff_0 ) : ( n394 ) ;
assign n396 =  ( n18 ) ? ( slice_stream_buff_0 ) : ( n395 ) ;
assign n397 =  ( n9 ) ? ( slice_stream_buff_0 ) : ( n396 ) ;
assign n398 =  ( n4 ) ? ( slice_stream_buff_0 ) : ( n397 ) ;
assign n399 =  ( n28 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n400 =  ( n35 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_1 ) ;
assign n401 =  ( n30 ) ? ( n399 ) : ( n400 ) ;
assign n402 =  ( n23 ) ? ( slice_stream_buff_1 ) : ( n401 ) ;
assign n403 =  ( n18 ) ? ( slice_stream_buff_1 ) : ( n402 ) ;
assign n404 =  ( n9 ) ? ( slice_stream_buff_1 ) : ( n403 ) ;
assign n405 =  ( n4 ) ? ( slice_stream_buff_1 ) : ( n404 ) ;
assign n406 =  ( n79 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n407 =  ( n28 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n408 =  ( n35 ) ? ( slice_stream_empty ) : ( slice_stream_empty ) ;
assign n409 =  ( n30 ) ? ( n407 ) : ( n408 ) ;
assign n410 =  ( n23 ) ? ( n406 ) : ( n409 ) ;
assign n411 =  ( n18 ) ? ( slice_stream_empty ) : ( n410 ) ;
assign n412 =  ( n9 ) ? ( slice_stream_empty ) : ( n411 ) ;
assign n413 =  ( n4 ) ? ( slice_stream_empty ) : ( n412 ) ;
assign n414 =  ( slice_stream_empty ) == ( 1'd1 )  ;
assign n415 =  ( n414 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n416 =  ( n28 ) ? ( 1'd0 ) : ( n415 ) ;
assign n417 =  ( n35 ) ? ( slice_stream_full ) : ( slice_stream_full ) ;
assign n418 =  ( n30 ) ? ( n416 ) : ( n417 ) ;
assign n419 =  ( n23 ) ? ( 1'd0 ) : ( n418 ) ;
assign n420 =  ( n18 ) ? ( slice_stream_full ) : ( n419 ) ;
assign n421 =  ( n9 ) ? ( slice_stream_full ) : ( n420 ) ;
assign n422 =  ( n4 ) ? ( slice_stream_full ) : ( n421 ) ;
assign n423 =  ( LB2D_shift_x ) >= ( 9'd8 )  ;
assign n424 = n80[71:64] ;
assign n425 = LB2D_shift_0[71:64] ;
assign n426 = LB2D_shift_1[71:64] ;
assign n427 = LB2D_shift_2[71:64] ;
assign n428 = LB2D_shift_3[71:64] ;
assign n429 = LB2D_shift_4[71:64] ;
assign n430 = LB2D_shift_5[71:64] ;
assign n431 = LB2D_shift_6[71:64] ;
assign n432 = LB2D_shift_7[71:64] ;
assign n433 =  { ( n431 ) , ( n432 ) }  ;
assign n434 =  { ( n430 ) , ( n433 ) }  ;
assign n435 =  { ( n429 ) , ( n434 ) }  ;
assign n436 =  { ( n428 ) , ( n435 ) }  ;
assign n437 =  { ( n427 ) , ( n436 ) }  ;
assign n438 =  { ( n426 ) , ( n437 ) }  ;
assign n439 =  { ( n425 ) , ( n438 ) }  ;
assign n440 =  { ( n424 ) , ( n439 ) }  ;
assign n441 = n80[63:56] ;
assign n442 = LB2D_shift_0[63:56] ;
assign n443 = LB2D_shift_1[63:56] ;
assign n444 = LB2D_shift_2[63:56] ;
assign n445 = LB2D_shift_3[63:56] ;
assign n446 = LB2D_shift_4[63:56] ;
assign n447 = LB2D_shift_5[63:56] ;
assign n448 = LB2D_shift_6[63:56] ;
assign n449 = LB2D_shift_7[63:56] ;
assign n450 =  { ( n448 ) , ( n449 ) }  ;
assign n451 =  { ( n447 ) , ( n450 ) }  ;
assign n452 =  { ( n446 ) , ( n451 ) }  ;
assign n453 =  { ( n445 ) , ( n452 ) }  ;
assign n454 =  { ( n444 ) , ( n453 ) }  ;
assign n455 =  { ( n443 ) , ( n454 ) }  ;
assign n456 =  { ( n442 ) , ( n455 ) }  ;
assign n457 =  { ( n441 ) , ( n456 ) }  ;
assign n458 = n80[55:48] ;
assign n459 = LB2D_shift_0[55:48] ;
assign n460 = LB2D_shift_1[55:48] ;
assign n461 = LB2D_shift_2[55:48] ;
assign n462 = LB2D_shift_3[55:48] ;
assign n463 = LB2D_shift_4[55:48] ;
assign n464 = LB2D_shift_5[55:48] ;
assign n465 = LB2D_shift_6[55:48] ;
assign n466 = LB2D_shift_7[55:48] ;
assign n467 =  { ( n465 ) , ( n466 ) }  ;
assign n468 =  { ( n464 ) , ( n467 ) }  ;
assign n469 =  { ( n463 ) , ( n468 ) }  ;
assign n470 =  { ( n462 ) , ( n469 ) }  ;
assign n471 =  { ( n461 ) , ( n470 ) }  ;
assign n472 =  { ( n460 ) , ( n471 ) }  ;
assign n473 =  { ( n459 ) , ( n472 ) }  ;
assign n474 =  { ( n458 ) , ( n473 ) }  ;
assign n475 = n80[47:40] ;
assign n476 = LB2D_shift_0[47:40] ;
assign n477 = LB2D_shift_1[47:40] ;
assign n478 = LB2D_shift_2[47:40] ;
assign n479 = LB2D_shift_3[47:40] ;
assign n480 = LB2D_shift_4[47:40] ;
assign n481 = LB2D_shift_5[47:40] ;
assign n482 = LB2D_shift_6[47:40] ;
assign n483 = LB2D_shift_7[47:40] ;
assign n484 =  { ( n482 ) , ( n483 ) }  ;
assign n485 =  { ( n481 ) , ( n484 ) }  ;
assign n486 =  { ( n480 ) , ( n485 ) }  ;
assign n487 =  { ( n479 ) , ( n486 ) }  ;
assign n488 =  { ( n478 ) , ( n487 ) }  ;
assign n489 =  { ( n477 ) , ( n488 ) }  ;
assign n490 =  { ( n476 ) , ( n489 ) }  ;
assign n491 =  { ( n475 ) , ( n490 ) }  ;
assign n492 = n80[39:32] ;
assign n493 = LB2D_shift_0[39:32] ;
assign n494 = LB2D_shift_1[39:32] ;
assign n495 = LB2D_shift_2[39:32] ;
assign n496 = LB2D_shift_3[39:32] ;
assign n497 = LB2D_shift_4[39:32] ;
assign n498 = LB2D_shift_5[39:32] ;
assign n499 = LB2D_shift_6[39:32] ;
assign n500 = LB2D_shift_7[39:32] ;
assign n501 =  { ( n499 ) , ( n500 ) }  ;
assign n502 =  { ( n498 ) , ( n501 ) }  ;
assign n503 =  { ( n497 ) , ( n502 ) }  ;
assign n504 =  { ( n496 ) , ( n503 ) }  ;
assign n505 =  { ( n495 ) , ( n504 ) }  ;
assign n506 =  { ( n494 ) , ( n505 ) }  ;
assign n507 =  { ( n493 ) , ( n506 ) }  ;
assign n508 =  { ( n492 ) , ( n507 ) }  ;
assign n509 = n80[31:24] ;
assign n510 = LB2D_shift_0[31:24] ;
assign n511 = LB2D_shift_1[31:24] ;
assign n512 = LB2D_shift_2[31:24] ;
assign n513 = LB2D_shift_3[31:24] ;
assign n514 = LB2D_shift_4[31:24] ;
assign n515 = LB2D_shift_5[31:24] ;
assign n516 = LB2D_shift_6[31:24] ;
assign n517 = LB2D_shift_7[31:24] ;
assign n518 =  { ( n516 ) , ( n517 ) }  ;
assign n519 =  { ( n515 ) , ( n518 ) }  ;
assign n520 =  { ( n514 ) , ( n519 ) }  ;
assign n521 =  { ( n513 ) , ( n520 ) }  ;
assign n522 =  { ( n512 ) , ( n521 ) }  ;
assign n523 =  { ( n511 ) , ( n522 ) }  ;
assign n524 =  { ( n510 ) , ( n523 ) }  ;
assign n525 =  { ( n509 ) , ( n524 ) }  ;
assign n526 = n80[23:16] ;
assign n527 = LB2D_shift_0[23:16] ;
assign n528 = LB2D_shift_1[23:16] ;
assign n529 = LB2D_shift_2[23:16] ;
assign n530 = LB2D_shift_3[23:16] ;
assign n531 = LB2D_shift_4[23:16] ;
assign n532 = LB2D_shift_5[23:16] ;
assign n533 = LB2D_shift_6[23:16] ;
assign n534 = LB2D_shift_7[23:16] ;
assign n535 =  { ( n533 ) , ( n534 ) }  ;
assign n536 =  { ( n532 ) , ( n535 ) }  ;
assign n537 =  { ( n531 ) , ( n536 ) }  ;
assign n538 =  { ( n530 ) , ( n537 ) }  ;
assign n539 =  { ( n529 ) , ( n538 ) }  ;
assign n540 =  { ( n528 ) , ( n539 ) }  ;
assign n541 =  { ( n527 ) , ( n540 ) }  ;
assign n542 =  { ( n526 ) , ( n541 ) }  ;
assign n543 = n80[15:8] ;
assign n544 = LB2D_shift_0[15:8] ;
assign n545 = LB2D_shift_1[15:8] ;
assign n546 = LB2D_shift_2[15:8] ;
assign n547 = LB2D_shift_3[15:8] ;
assign n548 = LB2D_shift_4[15:8] ;
assign n549 = LB2D_shift_5[15:8] ;
assign n550 = LB2D_shift_6[15:8] ;
assign n551 = LB2D_shift_7[15:8] ;
assign n552 =  { ( n550 ) , ( n551 ) }  ;
assign n553 =  { ( n549 ) , ( n552 ) }  ;
assign n554 =  { ( n548 ) , ( n553 ) }  ;
assign n555 =  { ( n547 ) , ( n554 ) }  ;
assign n556 =  { ( n546 ) , ( n555 ) }  ;
assign n557 =  { ( n545 ) , ( n556 ) }  ;
assign n558 =  { ( n544 ) , ( n557 ) }  ;
assign n559 =  { ( n543 ) , ( n558 ) }  ;
assign n560 = n80[7:0] ;
assign n561 = LB2D_shift_0[7:0] ;
assign n562 = LB2D_shift_1[7:0] ;
assign n563 = LB2D_shift_2[7:0] ;
assign n564 = LB2D_shift_3[7:0] ;
assign n565 = LB2D_shift_4[7:0] ;
assign n566 = LB2D_shift_5[7:0] ;
assign n567 = LB2D_shift_6[7:0] ;
assign n568 = LB2D_shift_7[7:0] ;
assign n569 =  { ( n567 ) , ( n568 ) }  ;
assign n570 =  { ( n566 ) , ( n569 ) }  ;
assign n571 =  { ( n565 ) , ( n570 ) }  ;
assign n572 =  { ( n564 ) , ( n571 ) }  ;
assign n573 =  { ( n563 ) , ( n572 ) }  ;
assign n574 =  { ( n562 ) , ( n573 ) }  ;
assign n575 =  { ( n561 ) , ( n574 ) }  ;
assign n576 =  { ( n560 ) , ( n575 ) }  ;
assign n577 =  { ( n559 ) , ( n576 ) }  ;
assign n578 =  { ( n542 ) , ( n577 ) }  ;
assign n579 =  { ( n525 ) , ( n578 ) }  ;
assign n580 =  { ( n508 ) , ( n579 ) }  ;
assign n581 =  { ( n491 ) , ( n580 ) }  ;
assign n582 =  { ( n474 ) , ( n581 ) }  ;
assign n583 =  { ( n457 ) , ( n582 ) }  ;
assign n584 =  { ( n440 ) , ( n583 ) }  ;
assign n585 =  ( n423 ) ? ( n584 ) : ( stencil_stream_buff_0 ) ;
assign n586 =  ( n35 ) ? ( stencil_stream_buff_0 ) : ( stencil_stream_buff_0 ) ;
assign n587 =  ( n30 ) ? ( stencil_stream_buff_0 ) : ( n586 ) ;
assign n588 =  ( n23 ) ? ( n585 ) : ( n587 ) ;
assign n589 =  ( n18 ) ? ( stencil_stream_buff_0 ) : ( n588 ) ;
assign n590 =  ( n9 ) ? ( stencil_stream_buff_0 ) : ( n589 ) ;
assign n591 =  ( n4 ) ? ( stencil_stream_buff_0 ) : ( n590 ) ;
assign n592 =  ( n35 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_1 ) ;
assign n593 =  ( n30 ) ? ( stencil_stream_buff_1 ) : ( n592 ) ;
assign n594 =  ( n23 ) ? ( stencil_stream_buff_0 ) : ( n593 ) ;
assign n595 =  ( n18 ) ? ( stencil_stream_buff_1 ) : ( n594 ) ;
assign n596 =  ( n9 ) ? ( stencil_stream_buff_1 ) : ( n595 ) ;
assign n597 =  ( n4 ) ? ( stencil_stream_buff_1 ) : ( n596 ) ;
assign n598 =  ( n148 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n599 =  ( n21 ) ? ( stencil_stream_empty ) : ( 1'd0 ) ;
assign n600 =  ( n35 ) ? ( stencil_stream_empty ) : ( stencil_stream_empty ) ;
assign n601 =  ( n30 ) ? ( stencil_stream_empty ) : ( n600 ) ;
assign n602 =  ( n23 ) ? ( n599 ) : ( n601 ) ;
assign n603 =  ( n18 ) ? ( n598 ) : ( n602 ) ;
assign n604 =  ( n9 ) ? ( stencil_stream_empty ) : ( n603 ) ;
assign n605 =  ( n4 ) ? ( stencil_stream_empty ) : ( n604 ) ;
assign n606 =  ( n14 ) ? ( 1'd0 ) : ( 1'd0 ) ;
assign n607 =  ( stencil_stream_empty ) == ( 1'd1 )  ;
assign n608 =  ( n607 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n609 =  ( n21 ) ? ( stencil_stream_full ) : ( n608 ) ;
assign n610 =  ( n35 ) ? ( stencil_stream_full ) : ( stencil_stream_full ) ;
assign n611 =  ( n30 ) ? ( stencil_stream_full ) : ( n610 ) ;
assign n612 =  ( n23 ) ? ( n609 ) : ( n611 ) ;
assign n613 =  ( n18 ) ? ( n606 ) : ( n612 ) ;
assign n614 =  ( n9 ) ? ( stencil_stream_full ) : ( n613 ) ;
assign n615 =  ( n4 ) ? ( stencil_stream_full ) : ( n614 ) ;
assign n616 = ~ ( n4 ) ;
assign n617 = ~ ( n9 ) ;
assign n618 =  ( n616 ) & ( n617 )  ;
assign n619 = ~ ( n18 ) ;
assign n620 =  ( n618 ) & ( n619 )  ;
assign n621 = ~ ( n23 ) ;
assign n622 =  ( n620 ) & ( n621 )  ;
assign n623 = ~ ( n30 ) ;
assign n624 =  ( n622 ) & ( n623 )  ;
assign n625 = ~ ( n35 ) ;
assign n626 =  ( n624 ) & ( n625 )  ;
assign n627 =  ( n624 ) & ( n35 )  ;
assign n628 =  ( n622 ) & ( n30 )  ;
assign n629 = ~ ( n313 ) ;
assign n630 =  ( n628 ) & ( n629 )  ;
assign n631 =  ( n628 ) & ( n313 )  ;
assign n632 =  ( n620 ) & ( n23 )  ;
assign n633 =  ( n618 ) & ( n18 )  ;
assign n634 =  ( n616 ) & ( n9 )  ;
assign LB2D_proc_0_addr0 = n631 ? (LB2D_proc_x) : (0);
assign LB2D_proc_0_data0 = n631 ? (n312) : (LB2D_proc_0[0]);
assign n635 = ~ ( n315 ) ;
assign n636 =  ( n628 ) & ( n635 )  ;
assign n637 =  ( n628 ) & ( n315 )  ;
assign LB2D_proc_1_addr0 = n637 ? (LB2D_proc_x) : (0);
assign LB2D_proc_1_data0 = n637 ? (n312) : (LB2D_proc_1[0]);
assign n638 = ~ ( n317 ) ;
assign n639 =  ( n628 ) & ( n638 )  ;
assign n640 =  ( n628 ) & ( n317 )  ;
assign LB2D_proc_2_addr0 = n640 ? (LB2D_proc_x) : (0);
assign LB2D_proc_2_data0 = n640 ? (n312) : (LB2D_proc_2[0]);
assign n641 = ~ ( n319 ) ;
assign n642 =  ( n628 ) & ( n641 )  ;
assign n643 =  ( n628 ) & ( n319 )  ;
assign LB2D_proc_3_addr0 = n643 ? (LB2D_proc_x) : (0);
assign LB2D_proc_3_data0 = n643 ? (n312) : (LB2D_proc_3[0]);
assign n644 = ~ ( n321 ) ;
assign n645 =  ( n628 ) & ( n644 )  ;
assign n646 =  ( n628 ) & ( n321 )  ;
assign LB2D_proc_4_addr0 = n646 ? (LB2D_proc_x) : (0);
assign LB2D_proc_4_data0 = n646 ? (n312) : (LB2D_proc_4[0]);
assign n647 = ~ ( n323 ) ;
assign n648 =  ( n628 ) & ( n647 )  ;
assign n649 =  ( n628 ) & ( n323 )  ;
assign LB2D_proc_5_addr0 = n649 ? (LB2D_proc_x) : (0);
assign LB2D_proc_5_data0 = n649 ? (n312) : (LB2D_proc_5[0]);
assign n650 = ~ ( n325 ) ;
assign n651 =  ( n628 ) & ( n650 )  ;
assign n652 =  ( n628 ) & ( n325 )  ;
assign LB2D_proc_6_addr0 = n652 ? (LB2D_proc_x) : (0);
assign LB2D_proc_6_data0 = n652 ? (n312) : (LB2D_proc_6[0]);
assign n653 =  ( LB2D_proc_w ) == ( 64'd7 )  ;
assign n654 = ~ ( n653 ) ;
assign n655 =  ( n628 ) & ( n654 )  ;
assign n656 =  ( n628 ) & ( n653 )  ;
assign LB2D_proc_7_addr0 = n656 ? (LB2D_proc_x) : (0);
assign LB2D_proc_7_data0 = n656 ? (n312) : (LB2D_proc_7[0]);
/*
function [7:0] gb_fun ;
input [647:0] arg0;
    begin
//TODO: Add the specific function HERE.    end
endfunction
*/

always @(posedge clk) begin
   if(rst) begin
       LB1D_buff <= LB1D_buff;
       LB1D_p_cnt <= LB1D_p_cnt;
       LB2D_proc_w <= LB2D_proc_w;
       LB2D_proc_x <= LB2D_proc_x;
       LB2D_proc_y <= LB2D_proc_y;
       LB2D_shift_0 <= LB2D_shift_0;
       LB2D_shift_1 <= LB2D_shift_1;
       LB2D_shift_2 <= LB2D_shift_2;
       LB2D_shift_3 <= LB2D_shift_3;
       LB2D_shift_4 <= LB2D_shift_4;
       LB2D_shift_5 <= LB2D_shift_5;
       LB2D_shift_6 <= LB2D_shift_6;
       LB2D_shift_7 <= LB2D_shift_7;
       LB2D_shift_x <= LB2D_shift_x;
       LB2D_shift_y <= LB2D_shift_y;
       arg_0_TDATA <= arg_0_TDATA;
       arg_0_TVALID <= arg_0_TVALID;
       arg_1_TREADY <= arg_1_TREADY;
       gb_exit_it_1 <= gb_exit_it_1;
       gb_exit_it_2 <= gb_exit_it_2;
       gb_exit_it_3 <= gb_exit_it_3;
       gb_exit_it_4 <= gb_exit_it_4;
       gb_exit_it_5 <= gb_exit_it_5;
       gb_exit_it_6 <= gb_exit_it_6;
       gb_exit_it_7 <= gb_exit_it_7;
       gb_exit_it_8 <= gb_exit_it_8;
       gb_p_cnt <= gb_p_cnt;
       gb_pp_it_1 <= gb_pp_it_1;
       gb_pp_it_2 <= gb_pp_it_2;
       gb_pp_it_3 <= gb_pp_it_3;
       gb_pp_it_4 <= gb_pp_it_4;
       gb_pp_it_5 <= gb_pp_it_5;
       gb_pp_it_6 <= gb_pp_it_6;
       gb_pp_it_7 <= gb_pp_it_7;
       gb_pp_it_8 <= gb_pp_it_8;
       gb_pp_it_9 <= gb_pp_it_9;
       in_stream_buff_0 <= in_stream_buff_0;
       in_stream_buff_1 <= in_stream_buff_1;
       in_stream_empty <= in_stream_empty;
       in_stream_full <= in_stream_full;
       slice_stream_buff_0 <= slice_stream_buff_0;
       slice_stream_buff_1 <= slice_stream_buff_1;
       slice_stream_empty <= slice_stream_empty;
       slice_stream_full <= slice_stream_full;
       stencil_stream_buff_0 <= stencil_stream_buff_0;
       stencil_stream_buff_1 <= stencil_stream_buff_1;
       stencil_stream_empty <= stencil_stream_empty;
       stencil_stream_full <= stencil_stream_full;
   end
   else if(step) begin
       LB1D_buff <= n41;
       LB1D_p_cnt <= n48;
       LB2D_proc_w <= n59;
       LB2D_proc_x <= n70;
       LB2D_proc_y <= n78;
       LB2D_shift_0 <= n86;
       LB2D_shift_1 <= n92;
       LB2D_shift_2 <= n98;
       LB2D_shift_3 <= n104;
       LB2D_shift_4 <= n110;
       LB2D_shift_5 <= n116;
       LB2D_shift_6 <= n122;
       LB2D_shift_7 <= n128;
       LB2D_shift_x <= n137;
       LB2D_shift_y <= n147;
       arg_0_TDATA <= n156;
       arg_0_TVALID <= n164;
       arg_1_TREADY <= n170;
       gb_exit_it_1 <= n179;
       gb_exit_it_2 <= n185;
       gb_exit_it_3 <= n191;
       gb_exit_it_4 <= n197;
       gb_exit_it_5 <= n203;
       gb_exit_it_6 <= n209;
       gb_exit_it_7 <= n215;
       gb_exit_it_8 <= n221;
       gb_p_cnt <= n229;
       gb_pp_it_1 <= n235;
       gb_pp_it_2 <= n241;
       gb_pp_it_3 <= n247;
       gb_pp_it_4 <= n253;
       gb_pp_it_5 <= n259;
       gb_pp_it_6 <= n265;
       gb_pp_it_7 <= n271;
       gb_pp_it_8 <= n277;
       gb_pp_it_9 <= n283;
       in_stream_buff_0 <= n289;
       in_stream_buff_1 <= n295;
       in_stream_empty <= n303;
       in_stream_full <= n311;
       slice_stream_buff_0 <= n398;
       slice_stream_buff_1 <= n405;
       slice_stream_empty <= n413;
       slice_stream_full <= n422;
       stencil_stream_buff_0 <= n591;
       stencil_stream_buff_1 <= n597;
       stencil_stream_empty <= n605;
       stencil_stream_full <= n615;
       LB2D_proc_0 [ LB2D_proc_0_addr0 ] <= LB2D_proc_0_data0;
       LB2D_proc_1 [ LB2D_proc_1_addr0 ] <= LB2D_proc_1_data0;
       LB2D_proc_2 [ LB2D_proc_2_addr0 ] <= LB2D_proc_2_data0;
       LB2D_proc_3 [ LB2D_proc_3_addr0 ] <= LB2D_proc_3_data0;
       LB2D_proc_4 [ LB2D_proc_4_addr0 ] <= LB2D_proc_4_data0;
       LB2D_proc_5 [ LB2D_proc_5_addr0 ] <= LB2D_proc_5_data0;
       LB2D_proc_6 [ LB2D_proc_6_addr0 ] <= LB2D_proc_6_data0;
       LB2D_proc_7 [ LB2D_proc_7_addr0 ] <= LB2D_proc_7_data0;
   end
end
endmodule
