module A(input clk, input rst, input in, output out);


endmodule

module B(input clk, input rst, input in, output out);


endmodule
