/* PREHEADER */
module fun_gb_fun (
    input [647:0] arg1,
    output [7:0] result
);
//TODO: Add the specific function HERE.
endmodule

/* END OF PREHEADER */
module SPEC_B(
arg_0_TREADY,
arg_1_TDATA,
arg_1_TVALID,
LB1D_buff,
LB1D_in,
LB1D_it_1,
LB1D_p_cnt,
LB1D_uIn,
LB2D_proc_w,
LB2D_proc_x,
LB2D_proc_y,
LB2D_shift_0,
LB2D_shift_1,
LB2D_shift_2,
LB2D_shift_3,
LB2D_shift_4,
LB2D_shift_5,
LB2D_shift_6,
LB2D_shift_7,
LB2D_shift_x,
LB2D_shift_y,
arg_0_TDATA,
arg_0_TVALID,
arg_1_TREADY,
gb_exit_it_1,
gb_exit_it_2,
gb_exit_it_3,
gb_exit_it_4,
gb_exit_it_5,
gb_exit_it_6,
gb_exit_it_7,
gb_exit_it_8,
gb_p_cnt,
gb_pp_it_1,
gb_pp_it_2,
gb_pp_it_3,
gb_pp_it_4,
gb_pp_it_5,
gb_pp_it_6,
gb_pp_it_7,
gb_pp_it_8,
gb_pp_it_9,
in_stream_buff_0,
in_stream_buff_1,
in_stream_empty,
in_stream_full,
slice_stream_buff_0,
slice_stream_buff_1,
slice_stream_empty,
slice_stream_full,
stencil_stream_buff_0,
stencil_stream_buff_1,
stencil_stream_empty,
stencil_stream_full,
clk,rst,
step
);
input            arg_0_TREADY;
input      [7:0] arg_1_TDATA;
input            arg_1_TVALID;
input clk;
input rst;
input step;
output      [7:0] LB1D_buff;
output      [7:0] LB1D_in;
output            LB1D_it_1;
output     [18:0] LB1D_p_cnt;
output      [7:0] LB1D_uIn;
output     [63:0] LB2D_proc_w;
output      [8:0] LB2D_proc_x;
output      [9:0] LB2D_proc_y;
output     [71:0] LB2D_shift_0;
output     [71:0] LB2D_shift_1;
output     [71:0] LB2D_shift_2;
output     [71:0] LB2D_shift_3;
output     [71:0] LB2D_shift_4;
output     [71:0] LB2D_shift_5;
output     [71:0] LB2D_shift_6;
output     [71:0] LB2D_shift_7;
output      [8:0] LB2D_shift_x;
output      [9:0] LB2D_shift_y;
output      [7:0] arg_0_TDATA;
output            arg_0_TVALID;
output            arg_1_TREADY;
output            gb_exit_it_1;
output            gb_exit_it_2;
output            gb_exit_it_3;
output            gb_exit_it_4;
output            gb_exit_it_5;
output            gb_exit_it_6;
output            gb_exit_it_7;
output            gb_exit_it_8;
output     [18:0] gb_p_cnt;
output            gb_pp_it_1;
output            gb_pp_it_2;
output            gb_pp_it_3;
output            gb_pp_it_4;
output            gb_pp_it_5;
output            gb_pp_it_6;
output            gb_pp_it_7;
output            gb_pp_it_8;
output            gb_pp_it_9;
output      [7:0] in_stream_buff_0;
output      [7:0] in_stream_buff_1;
output            in_stream_empty;
output            in_stream_full;
output     [71:0] slice_stream_buff_0;
output     [71:0] slice_stream_buff_1;
output            slice_stream_empty;
output            slice_stream_full;
output    [647:0] stencil_stream_buff_0;
output    [647:0] stencil_stream_buff_1;
output            stencil_stream_empty;
output            stencil_stream_full;
reg      [7:0] LB1D_buff;
reg      [7:0] LB1D_in;
reg            LB1D_it_1;
reg     [18:0] LB1D_p_cnt;
reg      [7:0] LB1D_uIn;
reg     [63:0] LB2D_proc_w;
reg      [8:0] LB2D_proc_x;
reg      [9:0] LB2D_proc_y;
reg     [71:0] LB2D_shift_0;
reg     [71:0] LB2D_shift_1;
reg     [71:0] LB2D_shift_2;
reg     [71:0] LB2D_shift_3;
reg     [71:0] LB2D_shift_4;
reg     [71:0] LB2D_shift_5;
reg     [71:0] LB2D_shift_6;
reg     [71:0] LB2D_shift_7;
reg      [8:0] LB2D_shift_x;
reg      [9:0] LB2D_shift_y;
reg      [7:0] arg_0_TDATA;
reg            arg_0_TVALID;
reg            arg_1_TREADY;
reg            gb_exit_it_1;
reg            gb_exit_it_2;
reg            gb_exit_it_3;
reg            gb_exit_it_4;
reg            gb_exit_it_5;
reg            gb_exit_it_6;
reg            gb_exit_it_7;
reg            gb_exit_it_8;
reg     [18:0] gb_p_cnt;
reg            gb_pp_it_1;
reg            gb_pp_it_2;
reg            gb_pp_it_3;
reg            gb_pp_it_4;
reg            gb_pp_it_5;
reg            gb_pp_it_6;
reg            gb_pp_it_7;
reg            gb_pp_it_8;
reg            gb_pp_it_9;
reg      [7:0] in_stream_buff_0;
reg      [7:0] in_stream_buff_1;
reg            in_stream_empty;
reg            in_stream_full;
reg     [71:0] slice_stream_buff_0;
reg     [71:0] slice_stream_buff_1;
reg            slice_stream_empty;
reg            slice_stream_full;
reg    [647:0] stencil_stream_buff_0;
reg    [647:0] stencil_stream_buff_1;
reg            stencil_stream_empty;
reg            stencil_stream_full;
wire            arg_0_TREADY;
wire      [7:0] arg_1_TDATA;
wire            arg_1_TVALID;
wire            n0;
wire            n1;
wire            n2;
wire            n3;
wire            n4;
wire            n5;
wire            n6;
wire            n7;
wire            n8;
wire            n9;
wire            n10;
wire            n11;
wire            n12;
wire            n13;
wire            n14;
wire            n15;
wire            n16;
wire            n17;
wire            n18;
wire            n19;
wire            n20;
wire            n21;
wire            n22;
wire            n23;
wire            n24;
wire            n25;
wire            n26;
wire            n27;
wire            n28;
wire      [7:0] n29;
wire      [7:0] n30;
wire      [7:0] n31;
wire      [7:0] n32;
wire      [7:0] n33;
wire      [7:0] n34;
wire      [7:0] n35;
wire      [7:0] n36;
wire      [7:0] n37;
wire      [7:0] n38;
wire            n39;
wire            n40;
wire            n41;
wire            n42;
wire            n43;
wire     [18:0] n44;
wire     [18:0] n45;
wire     [18:0] n46;
wire     [18:0] n47;
wire     [18:0] n48;
wire     [18:0] n49;
wire     [18:0] n50;
wire      [7:0] n51;
wire      [7:0] n52;
wire      [7:0] n53;
wire      [7:0] n54;
wire            n55;
wire            n56;
wire     [63:0] n57;
wire     [63:0] n58;
wire     [63:0] n59;
wire     [63:0] n60;
wire     [63:0] n61;
wire     [63:0] n62;
wire     [63:0] n63;
wire     [63:0] n64;
wire      [8:0] n65;
wire      [8:0] n66;
wire      [8:0] n67;
wire      [8:0] n68;
wire      [8:0] n69;
wire      [8:0] n70;
wire      [8:0] n71;
wire            n72;
wire      [9:0] n73;
wire      [9:0] n74;
wire      [9:0] n75;
wire      [9:0] n76;
wire      [9:0] n77;
wire      [9:0] n78;
wire      [9:0] n79;
wire      [9:0] n80;
wire     [71:0] n81;
wire     [71:0] n82;
wire     [71:0] n83;
wire     [71:0] n84;
wire     [71:0] n85;
wire     [71:0] n86;
wire     [71:0] n87;
wire     [71:0] n88;
wire     [71:0] n89;
wire     [71:0] n90;
wire     [71:0] n91;
wire     [71:0] n92;
wire     [71:0] n93;
wire     [71:0] n94;
wire     [71:0] n95;
wire     [71:0] n96;
wire     [71:0] n97;
wire     [71:0] n98;
wire     [71:0] n99;
wire     [71:0] n100;
wire     [71:0] n101;
wire     [71:0] n102;
wire     [71:0] n103;
wire     [71:0] n104;
wire     [71:0] n105;
wire     [71:0] n106;
wire     [71:0] n107;
wire     [71:0] n108;
wire     [71:0] n109;
wire     [71:0] n110;
wire     [71:0] n111;
wire     [71:0] n112;
wire     [71:0] n113;
wire     [71:0] n114;
wire     [71:0] n115;
wire            n116;
wire     [71:0] n117;
wire     [71:0] n118;
wire     [71:0] n119;
wire     [71:0] n120;
wire     [71:0] n121;
wire     [71:0] n122;
wire            n123;
wire      [8:0] n124;
wire      [8:0] n125;
wire      [8:0] n126;
wire      [8:0] n127;
wire      [8:0] n128;
wire      [8:0] n129;
wire      [8:0] n130;
wire            n131;
wire            n132;
wire      [9:0] n133;
wire      [9:0] n134;
wire      [9:0] n135;
wire      [9:0] n136;
wire      [9:0] n137;
wire      [9:0] n138;
wire      [9:0] n139;
wire      [9:0] n140;
wire            n141;
wire    [647:0] n142;
wire      [7:0] n143;
wire      [7:0] n145;
wire      [7:0] n146;
wire      [7:0] n147;
wire      [7:0] n148;
wire      [7:0] n149;
wire      [7:0] n150;
wire            n151;
wire            n152;
wire            n153;
wire            n154;
wire            n155;
wire            n156;
wire            n157;
wire            n158;
wire            n159;
wire            n160;
wire            n161;
wire            n162;
wire            n163;
wire            n164;
wire            n165;
wire            n166;
wire            n167;
wire            n168;
wire            n169;
wire            n170;
wire            n171;
wire            n172;
wire            n173;
wire            n174;
wire            n175;
wire            n176;
wire            n177;
wire            n178;
wire            n179;
wire            n180;
wire            n181;
wire            n182;
wire            n183;
wire            n184;
wire            n185;
wire            n186;
wire            n187;
wire            n188;
wire            n189;
wire            n190;
wire            n191;
wire            n192;
wire            n193;
wire            n194;
wire            n195;
wire            n196;
wire            n197;
wire            n198;
wire            n199;
wire            n200;
wire            n201;
wire            n202;
wire            n203;
wire            n204;
wire            n205;
wire            n206;
wire            n207;
wire     [18:0] n208;
wire     [18:0] n209;
wire     [18:0] n210;
wire     [18:0] n211;
wire     [18:0] n212;
wire     [18:0] n213;
wire     [18:0] n214;
wire            n215;
wire            n216;
wire            n217;
wire            n218;
wire            n219;
wire            n220;
wire            n221;
wire            n222;
wire            n223;
wire            n224;
wire            n225;
wire            n226;
wire            n227;
wire            n228;
wire            n229;
wire            n230;
wire            n231;
wire            n232;
wire            n233;
wire            n234;
wire            n235;
wire            n236;
wire            n237;
wire            n238;
wire            n239;
wire            n240;
wire            n241;
wire            n242;
wire            n243;
wire            n244;
wire            n245;
wire            n246;
wire            n247;
wire            n248;
wire            n249;
wire            n250;
wire            n251;
wire            n252;
wire            n253;
wire            n254;
wire            n255;
wire            n256;
wire            n257;
wire            n258;
wire            n259;
wire      [7:0] n260;
wire      [7:0] n261;
wire      [7:0] n262;
wire      [7:0] n263;
wire      [7:0] n264;
wire      [7:0] n265;
wire      [7:0] n266;
wire      [7:0] n267;
wire      [7:0] n268;
wire      [7:0] n269;
wire            n270;
wire            n271;
wire            n272;
wire            n273;
wire            n274;
wire            n275;
wire            n276;
wire            n277;
wire            n278;
wire            n279;
wire            n280;
wire            n281;
wire            n282;
wire            n283;
wire      [7:0] n284;
wire            n285;
wire      [8:0] n286;
wire      [7:0] n287;
wire            n288;
wire      [7:0] n289;
wire            n290;
wire      [7:0] n291;
wire            n292;
wire      [7:0] n293;
wire            n294;
wire      [7:0] n295;
wire            n296;
wire      [7:0] n297;
wire            n298;
wire      [7:0] n299;
wire      [7:0] n300;
wire      [7:0] n301;
wire      [7:0] n302;
wire      [7:0] n303;
wire      [7:0] n304;
wire      [7:0] n305;
wire      [7:0] n306;
wire      [7:0] n307;
wire      [7:0] n308;
wire      [7:0] n309;
wire      [7:0] n310;
wire      [7:0] n311;
wire      [7:0] n312;
wire      [7:0] n313;
wire      [7:0] n314;
wire      [7:0] n315;
wire      [7:0] n316;
wire      [7:0] n317;
wire      [7:0] n318;
wire      [7:0] n319;
wire      [7:0] n320;
wire      [7:0] n321;
wire      [7:0] n322;
wire      [7:0] n323;
wire      [7:0] n324;
wire      [7:0] n325;
wire      [7:0] n326;
wire      [7:0] n327;
wire      [7:0] n328;
wire      [7:0] n329;
wire      [7:0] n330;
wire      [7:0] n331;
wire      [7:0] n332;
wire      [7:0] n333;
wire      [7:0] n334;
wire      [7:0] n335;
wire      [7:0] n336;
wire      [7:0] n337;
wire      [7:0] n338;
wire      [7:0] n339;
wire      [7:0] n340;
wire      [7:0] n341;
wire      [7:0] n342;
wire      [7:0] n343;
wire      [7:0] n344;
wire      [7:0] n345;
wire      [7:0] n346;
wire      [7:0] n347;
wire      [7:0] n348;
wire      [7:0] n349;
wire      [7:0] n350;
wire      [7:0] n351;
wire      [7:0] n352;
wire      [7:0] n353;
wire      [7:0] n354;
wire      [7:0] n355;
wire      [7:0] n356;
wire     [15:0] n357;
wire     [23:0] n358;
wire     [31:0] n359;
wire     [39:0] n360;
wire     [47:0] n361;
wire     [55:0] n362;
wire     [63:0] n363;
wire     [71:0] n364;
wire     [71:0] n365;
wire     [71:0] n366;
wire     [71:0] n367;
wire     [71:0] n368;
wire     [71:0] n369;
wire     [71:0] n370;
wire     [71:0] n371;
wire     [71:0] n372;
wire     [71:0] n373;
wire     [71:0] n374;
wire     [71:0] n375;
wire     [71:0] n376;
wire            n377;
wire            n378;
wire            n379;
wire            n380;
wire            n381;
wire            n382;
wire            n383;
wire            n384;
wire            n385;
wire            n386;
wire            n387;
wire            n388;
wire            n389;
wire            n390;
wire            n391;
wire            n392;
wire            n393;
wire            n394;
wire      [7:0] n395;
wire      [7:0] n396;
wire      [7:0] n397;
wire      [7:0] n398;
wire      [7:0] n399;
wire      [7:0] n400;
wire      [7:0] n401;
wire      [7:0] n402;
wire      [7:0] n403;
wire     [15:0] n404;
wire     [23:0] n405;
wire     [31:0] n406;
wire     [39:0] n407;
wire     [47:0] n408;
wire     [55:0] n409;
wire     [63:0] n410;
wire     [71:0] n411;
wire      [7:0] n412;
wire      [7:0] n413;
wire      [7:0] n414;
wire      [7:0] n415;
wire      [7:0] n416;
wire      [7:0] n417;
wire      [7:0] n418;
wire      [7:0] n419;
wire      [7:0] n420;
wire     [15:0] n421;
wire     [23:0] n422;
wire     [31:0] n423;
wire     [39:0] n424;
wire     [47:0] n425;
wire     [55:0] n426;
wire     [63:0] n427;
wire     [71:0] n428;
wire      [7:0] n429;
wire      [7:0] n430;
wire      [7:0] n431;
wire      [7:0] n432;
wire      [7:0] n433;
wire      [7:0] n434;
wire      [7:0] n435;
wire      [7:0] n436;
wire      [7:0] n437;
wire     [15:0] n438;
wire     [23:0] n439;
wire     [31:0] n440;
wire     [39:0] n441;
wire     [47:0] n442;
wire     [55:0] n443;
wire     [63:0] n444;
wire     [71:0] n445;
wire      [7:0] n446;
wire      [7:0] n447;
wire      [7:0] n448;
wire      [7:0] n449;
wire      [7:0] n450;
wire      [7:0] n451;
wire      [7:0] n452;
wire      [7:0] n453;
wire      [7:0] n454;
wire     [15:0] n455;
wire     [23:0] n456;
wire     [31:0] n457;
wire     [39:0] n458;
wire     [47:0] n459;
wire     [55:0] n460;
wire     [63:0] n461;
wire     [71:0] n462;
wire      [7:0] n463;
wire      [7:0] n464;
wire      [7:0] n465;
wire      [7:0] n466;
wire      [7:0] n467;
wire      [7:0] n468;
wire      [7:0] n469;
wire      [7:0] n470;
wire      [7:0] n471;
wire     [15:0] n472;
wire     [23:0] n473;
wire     [31:0] n474;
wire     [39:0] n475;
wire     [47:0] n476;
wire     [55:0] n477;
wire     [63:0] n478;
wire     [71:0] n479;
wire      [7:0] n480;
wire      [7:0] n481;
wire      [7:0] n482;
wire      [7:0] n483;
wire      [7:0] n484;
wire      [7:0] n485;
wire      [7:0] n486;
wire      [7:0] n487;
wire      [7:0] n488;
wire     [15:0] n489;
wire     [23:0] n490;
wire     [31:0] n491;
wire     [39:0] n492;
wire     [47:0] n493;
wire     [55:0] n494;
wire     [63:0] n495;
wire     [71:0] n496;
wire      [7:0] n497;
wire      [7:0] n498;
wire      [7:0] n499;
wire      [7:0] n500;
wire      [7:0] n501;
wire      [7:0] n502;
wire      [7:0] n503;
wire      [7:0] n504;
wire      [7:0] n505;
wire     [15:0] n506;
wire     [23:0] n507;
wire     [31:0] n508;
wire     [39:0] n509;
wire     [47:0] n510;
wire     [55:0] n511;
wire     [63:0] n512;
wire     [71:0] n513;
wire      [7:0] n514;
wire      [7:0] n515;
wire      [7:0] n516;
wire      [7:0] n517;
wire      [7:0] n518;
wire      [7:0] n519;
wire      [7:0] n520;
wire      [7:0] n521;
wire      [7:0] n522;
wire     [15:0] n523;
wire     [23:0] n524;
wire     [31:0] n525;
wire     [39:0] n526;
wire     [47:0] n527;
wire     [55:0] n528;
wire     [63:0] n529;
wire     [71:0] n530;
wire      [7:0] n531;
wire      [7:0] n532;
wire      [7:0] n533;
wire      [7:0] n534;
wire      [7:0] n535;
wire      [7:0] n536;
wire      [7:0] n537;
wire      [7:0] n538;
wire      [7:0] n539;
wire     [15:0] n540;
wire     [23:0] n541;
wire     [31:0] n542;
wire     [39:0] n543;
wire     [47:0] n544;
wire     [55:0] n545;
wire     [63:0] n546;
wire     [71:0] n547;
wire    [143:0] n548;
wire    [215:0] n549;
wire    [287:0] n550;
wire    [359:0] n551;
wire    [431:0] n552;
wire    [503:0] n553;
wire    [575:0] n554;
wire    [647:0] n555;
wire    [647:0] n556;
wire    [647:0] n557;
wire    [647:0] n558;
wire    [647:0] n559;
wire    [647:0] n560;
wire    [647:0] n561;
wire            n562;
wire    [647:0] n563;
wire    [647:0] n564;
wire    [647:0] n565;
wire    [647:0] n566;
wire    [647:0] n567;
wire            n568;
wire            n569;
wire            n570;
wire            n571;
wire            n572;
wire            n573;
wire            n574;
wire            n575;
wire            n576;
wire            n577;
wire            n578;
wire            n579;
wire            n580;
wire            n581;
wire            n582;
wire            n583;
wire            n584;
wire      [8:0] LB2D_proc_0_addr0;
wire      [7:0] LB2D_proc_0_data0;
wire            LB2D_proc_0_wen0;
wire            n585;
wire            n586;
wire            n587;
wire            n588;
wire            n589;
wire            n590;
wire            n591;
wire            n592;
wire            n593;
wire            n594;
wire            n595;
wire            n596;
wire            n597;
wire            n598;
wire            n599;
wire            n600;
wire            n601;
wire            n602;
wire      [8:0] LB2D_proc_1_addr0;
wire      [7:0] LB2D_proc_1_data0;
wire            LB2D_proc_1_wen0;
wire            n603;
wire            n604;
wire            n605;
wire      [8:0] LB2D_proc_2_addr0;
wire      [7:0] LB2D_proc_2_data0;
wire            LB2D_proc_2_wen0;
wire            n606;
wire            n607;
wire            n608;
wire      [8:0] LB2D_proc_3_addr0;
wire      [7:0] LB2D_proc_3_data0;
wire            LB2D_proc_3_wen0;
wire            n609;
wire            n610;
wire            n611;
wire      [8:0] LB2D_proc_4_addr0;
wire      [7:0] LB2D_proc_4_data0;
wire            LB2D_proc_4_wen0;
wire            n612;
wire            n613;
wire            n614;
wire      [8:0] LB2D_proc_5_addr0;
wire      [7:0] LB2D_proc_5_data0;
wire            LB2D_proc_5_wen0;
wire            n615;
wire            n616;
wire            n617;
wire      [8:0] LB2D_proc_6_addr0;
wire      [7:0] LB2D_proc_6_data0;
wire            LB2D_proc_6_wen0;
wire            n618;
wire            n619;
wire            n620;
wire      [8:0] LB2D_proc_7_addr0;
wire      [7:0] LB2D_proc_7_data0;
wire            LB2D_proc_7_wen0;
wire            n621;
wire            n622;
wire            n623;
reg      [7:0] LB2D_proc_0[511:0];
reg      [7:0] LB2D_proc_1[511:0];
reg      [7:0] LB2D_proc_2[511:0];
reg      [7:0] LB2D_proc_3[511:0];
reg      [7:0] LB2D_proc_4[511:0];
reg      [7:0] LB2D_proc_5[511:0];
reg      [7:0] LB2D_proc_6[511:0];
reg      [7:0] LB2D_proc_7[511:0];
wire clk;
wire rst;
wire step;
assign n0 =  ( arg_0_TREADY ) == ( 1'd1 )  ;
assign n1 =  ( arg_0_TVALID ) == ( 1'd1 )  ;
assign n2 =  ( n0 ) & ( n1 )  ;
assign n3 =  ( arg_1_TVALID ) == ( 1'd0 )  ;
assign n4 =  ( n2 ) & ( n3 )  ;
assign n5 =  ( arg_0_TVALID ) == ( 1'd0 )  ;
assign n6 =  ( gb_exit_it_1 ) == ( 1'd0 )  ;
assign n7 =  ( stencil_stream_empty ) == ( 1'd0 )  ;
assign n8 =  ( n6 ) & ( n7 )  ;
assign n9 =  ( gb_exit_it_1 ) == ( 1'd1 )  ;
assign n10 =  ( gb_exit_it_8 ) == ( 1'd0 )  ;
assign n11 =  ( n9 ) & ( n10 )  ;
assign n12 =  ( n8 ) | ( n11 )  ;
assign n13 =  ( n5 ) & ( n12 )  ;
assign n14 =  ( slice_stream_empty ) == ( 1'd0 )  ;
assign n15 =  ( stencil_stream_full ) == ( 1'd0 )  ;
assign n16 =  ( LB2D_shift_x ) < ( 9'd8 )  ;
assign n17 =  ( LB2D_shift_x ) > ( 9'd0 )  ;
assign n18 =  ( n16 ) & ( n17 )  ;
assign n19 =  ( n15 ) | ( n18 )  ;
assign n20 =  ( n14 ) & ( n19 )  ;
assign n21 =  ( in_stream_empty ) == ( 1'd0 )  ;
assign n22 =  ( slice_stream_full ) == ( 1'd0 )  ;
assign n23 =  ( LB2D_proc_y ) < ( 10'd8 )  ;
assign n24 =  ( n22 ) | ( n23 )  ;
assign n25 =  ( n21 ) & ( n24 )  ;
assign n26 =  ( arg_1_TREADY ) == ( 1'd0 )  ;
assign n27 =  ( in_stream_full ) == ( 1'd0 )  ;
assign n28 =  ( n26 ) & ( n27 )  ;
assign n29 =  ( n28 ) ? ( LB1D_uIn ) : ( LB1D_buff ) ;
assign n30 =  ( n25 ) ? ( LB1D_buff ) : ( n29 ) ;
assign n31 =  ( n20 ) ? ( LB1D_buff ) : ( n30 ) ;
assign n32 =  ( n13 ) ? ( LB1D_buff ) : ( n31 ) ;
assign n33 =  ( n4 ) ? ( LB1D_buff ) : ( n32 ) ;
assign n34 =  ( n28 ) ? ( LB1D_in ) : ( LB1D_in ) ;
assign n35 =  ( n25 ) ? ( LB1D_in ) : ( n34 ) ;
assign n36 =  ( n20 ) ? ( LB1D_in ) : ( n35 ) ;
assign n37 =  ( n13 ) ? ( LB1D_in ) : ( n36 ) ;
assign n38 =  ( n4 ) ? ( LB1D_in ) : ( n37 ) ;
assign n39 =  ( LB1D_it_1 ) == ( 1'd1 )  ;
assign n40 =  ( LB1D_p_cnt ) == ( 19'd316224 )  ;
assign n41 =  ( n39 ) & ( n40 )  ;
assign n42 =  ( n41 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n43 =  ( n28 ) ? ( n42 ) : ( LB1D_it_1 ) ;
assign n44 =  ( LB1D_p_cnt ) + ( 19'd1 )  ;
assign n45 =  ( n41 ) ? ( 19'd0 ) : ( n44 ) ;
assign n46 =  ( n28 ) ? ( n45 ) : ( LB1D_p_cnt ) ;
assign n47 =  ( n25 ) ? ( LB1D_p_cnt ) : ( n46 ) ;
assign n48 =  ( n20 ) ? ( LB1D_p_cnt ) : ( n47 ) ;
assign n49 =  ( n13 ) ? ( LB1D_p_cnt ) : ( n48 ) ;
assign n50 =  ( n4 ) ? ( LB1D_p_cnt ) : ( n49 ) ;
assign n51 =  ( n28 ) ? ( LB1D_in ) : ( LB1D_uIn ) ;
assign n52 =  ( n25 ) ? ( LB1D_uIn ) : ( n51 ) ;
assign n53 =  ( n20 ) ? ( LB1D_uIn ) : ( n52 ) ;
assign n54 =  ( n13 ) ? ( LB1D_uIn ) : ( n53 ) ;
assign n55 =  ( LB2D_proc_x ) == ( 9'd488 )  ;
assign n56 =  ( LB2D_proc_w ) == ( 64'd7 )  ;
assign n57 =  ( LB2D_proc_w ) + ( 64'd1 )  ;
assign n58 =  ( n56 ) ? ( 64'd0 ) : ( n57 ) ;
assign n59 =  ( n55 ) ? ( n58 ) : ( LB2D_proc_w ) ;
assign n60 =  ( n28 ) ? ( LB2D_proc_w ) : ( LB2D_proc_w ) ;
assign n61 =  ( n25 ) ? ( n59 ) : ( n60 ) ;
assign n62 =  ( n20 ) ? ( LB2D_proc_w ) : ( n61 ) ;
assign n63 =  ( n13 ) ? ( LB2D_proc_w ) : ( n62 ) ;
assign n64 =  ( n4 ) ? ( LB2D_proc_w ) : ( n63 ) ;
assign n65 =  ( LB2D_proc_x ) + ( 9'd1 )  ;
assign n66 =  ( n55 ) ? ( 9'd1 ) : ( n65 ) ;
assign n67 =  ( n28 ) ? ( LB2D_proc_x ) : ( LB2D_proc_x ) ;
assign n68 =  ( n25 ) ? ( n66 ) : ( n67 ) ;
assign n69 =  ( n20 ) ? ( LB2D_proc_x ) : ( n68 ) ;
assign n70 =  ( n13 ) ? ( LB2D_proc_x ) : ( n69 ) ;
assign n71 =  ( n4 ) ? ( LB2D_proc_x ) : ( n70 ) ;
assign n72 =  ( LB2D_proc_y ) == ( 10'd648 )  ;
assign n73 =  ( LB2D_proc_y ) + ( 10'd1 )  ;
assign n74 =  ( n72 ) ? ( 10'd0 ) : ( n73 ) ;
assign n75 =  ( n55 ) ? ( n74 ) : ( LB2D_proc_y ) ;
assign n76 =  ( n28 ) ? ( LB2D_proc_y ) : ( LB2D_proc_y ) ;
assign n77 =  ( n25 ) ? ( n75 ) : ( n76 ) ;
assign n78 =  ( n20 ) ? ( LB2D_proc_y ) : ( n77 ) ;
assign n79 =  ( n13 ) ? ( LB2D_proc_y ) : ( n78 ) ;
assign n80 =  ( n4 ) ? ( LB2D_proc_y ) : ( n79 ) ;
assign n81 =  ( n28 ) ? ( LB2D_shift_0 ) : ( LB2D_shift_0 ) ;
assign n82 =  ( n25 ) ? ( LB2D_shift_0 ) : ( n81 ) ;
assign n83 =  ( n20 ) ? ( LB2D_shift_1 ) : ( n82 ) ;
assign n84 =  ( n13 ) ? ( LB2D_shift_0 ) : ( n83 ) ;
assign n85 =  ( n4 ) ? ( LB2D_shift_0 ) : ( n84 ) ;
assign n86 =  ( n28 ) ? ( LB2D_shift_1 ) : ( LB2D_shift_1 ) ;
assign n87 =  ( n25 ) ? ( LB2D_shift_1 ) : ( n86 ) ;
assign n88 =  ( n20 ) ? ( LB2D_shift_2 ) : ( n87 ) ;
assign n89 =  ( n13 ) ? ( LB2D_shift_1 ) : ( n88 ) ;
assign n90 =  ( n4 ) ? ( LB2D_shift_1 ) : ( n89 ) ;
assign n91 =  ( n28 ) ? ( LB2D_shift_2 ) : ( LB2D_shift_2 ) ;
assign n92 =  ( n25 ) ? ( LB2D_shift_2 ) : ( n91 ) ;
assign n93 =  ( n20 ) ? ( LB2D_shift_3 ) : ( n92 ) ;
assign n94 =  ( n13 ) ? ( LB2D_shift_2 ) : ( n93 ) ;
assign n95 =  ( n4 ) ? ( LB2D_shift_2 ) : ( n94 ) ;
assign n96 =  ( n28 ) ? ( LB2D_shift_3 ) : ( LB2D_shift_3 ) ;
assign n97 =  ( n25 ) ? ( LB2D_shift_3 ) : ( n96 ) ;
assign n98 =  ( n20 ) ? ( LB2D_shift_4 ) : ( n97 ) ;
assign n99 =  ( n13 ) ? ( LB2D_shift_3 ) : ( n98 ) ;
assign n100 =  ( n4 ) ? ( LB2D_shift_3 ) : ( n99 ) ;
assign n101 =  ( n28 ) ? ( LB2D_shift_4 ) : ( LB2D_shift_4 ) ;
assign n102 =  ( n25 ) ? ( LB2D_shift_4 ) : ( n101 ) ;
assign n103 =  ( n20 ) ? ( LB2D_shift_5 ) : ( n102 ) ;
assign n104 =  ( n13 ) ? ( LB2D_shift_4 ) : ( n103 ) ;
assign n105 =  ( n4 ) ? ( LB2D_shift_4 ) : ( n104 ) ;
assign n106 =  ( n28 ) ? ( LB2D_shift_5 ) : ( LB2D_shift_5 ) ;
assign n107 =  ( n25 ) ? ( LB2D_shift_5 ) : ( n106 ) ;
assign n108 =  ( n20 ) ? ( LB2D_shift_6 ) : ( n107 ) ;
assign n109 =  ( n13 ) ? ( LB2D_shift_5 ) : ( n108 ) ;
assign n110 =  ( n4 ) ? ( LB2D_shift_5 ) : ( n109 ) ;
assign n111 =  ( n28 ) ? ( LB2D_shift_6 ) : ( LB2D_shift_6 ) ;
assign n112 =  ( n25 ) ? ( LB2D_shift_6 ) : ( n111 ) ;
assign n113 =  ( n20 ) ? ( LB2D_shift_7 ) : ( n112 ) ;
assign n114 =  ( n13 ) ? ( LB2D_shift_6 ) : ( n113 ) ;
assign n115 =  ( n4 ) ? ( LB2D_shift_6 ) : ( n114 ) ;
assign n116 =  ( slice_stream_full ) == ( 1'd1 )  ;
assign n117 =  ( n116 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n118 =  ( n28 ) ? ( LB2D_shift_7 ) : ( LB2D_shift_7 ) ;
assign n119 =  ( n25 ) ? ( LB2D_shift_7 ) : ( n118 ) ;
assign n120 =  ( n20 ) ? ( n117 ) : ( n119 ) ;
assign n121 =  ( n13 ) ? ( LB2D_shift_7 ) : ( n120 ) ;
assign n122 =  ( n4 ) ? ( LB2D_shift_7 ) : ( n121 ) ;
assign n123 =  ( LB2D_shift_x ) == ( 9'd488 )  ;
assign n124 =  ( LB2D_shift_x ) + ( 9'd1 )  ;
assign n125 =  ( n123 ) ? ( 9'd0 ) : ( n124 ) ;
assign n126 =  ( n28 ) ? ( LB2D_shift_x ) : ( LB2D_shift_x ) ;
assign n127 =  ( n25 ) ? ( LB2D_shift_x ) : ( n126 ) ;
assign n128 =  ( n20 ) ? ( n125 ) : ( n127 ) ;
assign n129 =  ( n13 ) ? ( LB2D_shift_x ) : ( n128 ) ;
assign n130 =  ( n4 ) ? ( LB2D_shift_x ) : ( n129 ) ;
assign n131 =  ( LB2D_shift_y ) < ( 10'd640 )  ;
assign n132 =  ( LB2D_shift_x ) < ( 9'd488 )  ;
assign n133 =  ( LB2D_shift_y ) + ( 10'd1 )  ;
assign n134 =  ( n132 ) ? ( LB2D_shift_y ) : ( n133 ) ;
assign n135 =  ( n131 ) ? ( n134 ) : ( 10'd640 ) ;
assign n136 =  ( n28 ) ? ( LB2D_shift_y ) : ( LB2D_shift_y ) ;
assign n137 =  ( n25 ) ? ( LB2D_shift_y ) : ( n136 ) ;
assign n138 =  ( n20 ) ? ( n135 ) : ( n137 ) ;
assign n139 =  ( n13 ) ? ( LB2D_shift_y ) : ( n138 ) ;
assign n140 =  ( n4 ) ? ( LB2D_shift_y ) : ( n139 ) ;
assign n141 =  ( stencil_stream_full ) == ( 1'd1 )  ;
assign n142 =  ( n141 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_0 ) ;
fun_gb_fun  applyFunc_n144(
    .arg1( n142 ),
    .result( n143 )
);
assign n145 = n143 ;
assign n146 =  ( n28 ) ? ( arg_0_TDATA ) : ( arg_0_TDATA ) ;
assign n147 =  ( n25 ) ? ( arg_0_TDATA ) : ( n146 ) ;
assign n148 =  ( n20 ) ? ( arg_0_TDATA ) : ( n147 ) ;
assign n149 =  ( n13 ) ? ( n145 ) : ( n148 ) ;
assign n150 =  ( n4 ) ? ( arg_0_TDATA ) : ( n149 ) ;
assign n151 =  ( gb_pp_it_8 ) == ( 1'd1 )  ;
assign n152 =  ( gb_exit_it_7 ) == ( 1'd0 )  ;
assign n153 =  ( n151 ) & ( n152 )  ;
assign n154 =  ( n153 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n155 =  ( n28 ) ? ( arg_0_TVALID ) : ( arg_0_TVALID ) ;
assign n156 =  ( n25 ) ? ( arg_0_TVALID ) : ( n155 ) ;
assign n157 =  ( n20 ) ? ( arg_0_TVALID ) : ( n156 ) ;
assign n158 =  ( n13 ) ? ( n154 ) : ( n157 ) ;
assign n159 =  ( n4 ) ? ( 1'd0 ) : ( n158 ) ;
assign n160 =  ( n28 ) ? ( 1'd1 ) : ( arg_1_TREADY ) ;
assign n161 =  ( n25 ) ? ( arg_1_TREADY ) : ( n160 ) ;
assign n162 =  ( n20 ) ? ( arg_1_TREADY ) : ( n161 ) ;
assign n163 =  ( n13 ) ? ( arg_1_TREADY ) : ( n162 ) ;
assign n164 =  ( n4 ) ? ( arg_1_TREADY ) : ( n163 ) ;
assign n165 =  ( gb_p_cnt ) == ( 19'd307200 )  ;
assign n166 =  ( n165 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n167 =  ( n28 ) ? ( gb_exit_it_1 ) : ( gb_exit_it_1 ) ;
assign n168 =  ( n25 ) ? ( gb_exit_it_1 ) : ( n167 ) ;
assign n169 =  ( n20 ) ? ( gb_exit_it_1 ) : ( n168 ) ;
assign n170 =  ( n13 ) ? ( n166 ) : ( n169 ) ;
assign n171 =  ( n4 ) ? ( gb_exit_it_1 ) : ( n170 ) ;
assign n172 =  ( n28 ) ? ( gb_exit_it_2 ) : ( gb_exit_it_2 ) ;
assign n173 =  ( n25 ) ? ( gb_exit_it_2 ) : ( n172 ) ;
assign n174 =  ( n20 ) ? ( gb_exit_it_2 ) : ( n173 ) ;
assign n175 =  ( n13 ) ? ( gb_exit_it_1 ) : ( n174 ) ;
assign n176 =  ( n4 ) ? ( gb_exit_it_2 ) : ( n175 ) ;
assign n177 =  ( n28 ) ? ( gb_exit_it_3 ) : ( gb_exit_it_3 ) ;
assign n178 =  ( n25 ) ? ( gb_exit_it_3 ) : ( n177 ) ;
assign n179 =  ( n20 ) ? ( gb_exit_it_3 ) : ( n178 ) ;
assign n180 =  ( n13 ) ? ( gb_exit_it_2 ) : ( n179 ) ;
assign n181 =  ( n4 ) ? ( gb_exit_it_3 ) : ( n180 ) ;
assign n182 =  ( n28 ) ? ( gb_exit_it_4 ) : ( gb_exit_it_4 ) ;
assign n183 =  ( n25 ) ? ( gb_exit_it_4 ) : ( n182 ) ;
assign n184 =  ( n20 ) ? ( gb_exit_it_4 ) : ( n183 ) ;
assign n185 =  ( n13 ) ? ( gb_exit_it_3 ) : ( n184 ) ;
assign n186 =  ( n4 ) ? ( gb_exit_it_4 ) : ( n185 ) ;
assign n187 =  ( n28 ) ? ( gb_exit_it_5 ) : ( gb_exit_it_5 ) ;
assign n188 =  ( n25 ) ? ( gb_exit_it_5 ) : ( n187 ) ;
assign n189 =  ( n20 ) ? ( gb_exit_it_5 ) : ( n188 ) ;
assign n190 =  ( n13 ) ? ( gb_exit_it_4 ) : ( n189 ) ;
assign n191 =  ( n4 ) ? ( gb_exit_it_5 ) : ( n190 ) ;
assign n192 =  ( n28 ) ? ( gb_exit_it_6 ) : ( gb_exit_it_6 ) ;
assign n193 =  ( n25 ) ? ( gb_exit_it_6 ) : ( n192 ) ;
assign n194 =  ( n20 ) ? ( gb_exit_it_6 ) : ( n193 ) ;
assign n195 =  ( n13 ) ? ( gb_exit_it_5 ) : ( n194 ) ;
assign n196 =  ( n4 ) ? ( gb_exit_it_6 ) : ( n195 ) ;
assign n197 =  ( n28 ) ? ( gb_exit_it_7 ) : ( gb_exit_it_7 ) ;
assign n198 =  ( n25 ) ? ( gb_exit_it_7 ) : ( n197 ) ;
assign n199 =  ( n20 ) ? ( gb_exit_it_7 ) : ( n198 ) ;
assign n200 =  ( n13 ) ? ( gb_exit_it_6 ) : ( n199 ) ;
assign n201 =  ( n4 ) ? ( gb_exit_it_7 ) : ( n200 ) ;
assign n202 =  ( n28 ) ? ( gb_exit_it_8 ) : ( gb_exit_it_8 ) ;
assign n203 =  ( n25 ) ? ( gb_exit_it_8 ) : ( n202 ) ;
assign n204 =  ( n20 ) ? ( gb_exit_it_8 ) : ( n203 ) ;
assign n205 =  ( n13 ) ? ( gb_exit_it_7 ) : ( n204 ) ;
assign n206 =  ( n4 ) ? ( gb_exit_it_8 ) : ( n205 ) ;
assign n207 =  ( gb_p_cnt ) < ( 19'd307200 )  ;
assign n208 =  ( gb_p_cnt ) + ( 19'd1 )  ;
assign n209 =  ( n207 ) ? ( n208 ) : ( 19'd307200 ) ;
assign n210 =  ( n28 ) ? ( gb_p_cnt ) : ( gb_p_cnt ) ;
assign n211 =  ( n25 ) ? ( gb_p_cnt ) : ( n210 ) ;
assign n212 =  ( n20 ) ? ( gb_p_cnt ) : ( n211 ) ;
assign n213 =  ( n13 ) ? ( n209 ) : ( n212 ) ;
assign n214 =  ( n4 ) ? ( gb_p_cnt ) : ( n213 ) ;
assign n215 =  ( n28 ) ? ( gb_pp_it_1 ) : ( gb_pp_it_1 ) ;
assign n216 =  ( n25 ) ? ( gb_pp_it_1 ) : ( n215 ) ;
assign n217 =  ( n20 ) ? ( gb_pp_it_1 ) : ( n216 ) ;
assign n218 =  ( n13 ) ? ( 1'd1 ) : ( n217 ) ;
assign n219 =  ( n4 ) ? ( gb_pp_it_1 ) : ( n218 ) ;
assign n220 =  ( n28 ) ? ( gb_pp_it_2 ) : ( gb_pp_it_2 ) ;
assign n221 =  ( n25 ) ? ( gb_pp_it_2 ) : ( n220 ) ;
assign n222 =  ( n20 ) ? ( gb_pp_it_2 ) : ( n221 ) ;
assign n223 =  ( n13 ) ? ( gb_pp_it_1 ) : ( n222 ) ;
assign n224 =  ( n4 ) ? ( gb_pp_it_2 ) : ( n223 ) ;
assign n225 =  ( n28 ) ? ( gb_pp_it_3 ) : ( gb_pp_it_3 ) ;
assign n226 =  ( n25 ) ? ( gb_pp_it_3 ) : ( n225 ) ;
assign n227 =  ( n20 ) ? ( gb_pp_it_3 ) : ( n226 ) ;
assign n228 =  ( n13 ) ? ( gb_pp_it_2 ) : ( n227 ) ;
assign n229 =  ( n4 ) ? ( gb_pp_it_3 ) : ( n228 ) ;
assign n230 =  ( n28 ) ? ( gb_pp_it_4 ) : ( gb_pp_it_4 ) ;
assign n231 =  ( n25 ) ? ( gb_pp_it_4 ) : ( n230 ) ;
assign n232 =  ( n20 ) ? ( gb_pp_it_4 ) : ( n231 ) ;
assign n233 =  ( n13 ) ? ( gb_pp_it_3 ) : ( n232 ) ;
assign n234 =  ( n4 ) ? ( gb_pp_it_4 ) : ( n233 ) ;
assign n235 =  ( n28 ) ? ( gb_pp_it_5 ) : ( gb_pp_it_5 ) ;
assign n236 =  ( n25 ) ? ( gb_pp_it_5 ) : ( n235 ) ;
assign n237 =  ( n20 ) ? ( gb_pp_it_5 ) : ( n236 ) ;
assign n238 =  ( n13 ) ? ( gb_pp_it_4 ) : ( n237 ) ;
assign n239 =  ( n4 ) ? ( gb_pp_it_5 ) : ( n238 ) ;
assign n240 =  ( n28 ) ? ( gb_pp_it_6 ) : ( gb_pp_it_6 ) ;
assign n241 =  ( n25 ) ? ( gb_pp_it_6 ) : ( n240 ) ;
assign n242 =  ( n20 ) ? ( gb_pp_it_6 ) : ( n241 ) ;
assign n243 =  ( n13 ) ? ( gb_pp_it_5 ) : ( n242 ) ;
assign n244 =  ( n4 ) ? ( gb_pp_it_6 ) : ( n243 ) ;
assign n245 =  ( n28 ) ? ( gb_pp_it_7 ) : ( gb_pp_it_7 ) ;
assign n246 =  ( n25 ) ? ( gb_pp_it_7 ) : ( n245 ) ;
assign n247 =  ( n20 ) ? ( gb_pp_it_7 ) : ( n246 ) ;
assign n248 =  ( n13 ) ? ( gb_pp_it_6 ) : ( n247 ) ;
assign n249 =  ( n4 ) ? ( gb_pp_it_7 ) : ( n248 ) ;
assign n250 =  ( n28 ) ? ( gb_pp_it_8 ) : ( gb_pp_it_8 ) ;
assign n251 =  ( n25 ) ? ( gb_pp_it_8 ) : ( n250 ) ;
assign n252 =  ( n20 ) ? ( gb_pp_it_8 ) : ( n251 ) ;
assign n253 =  ( n13 ) ? ( gb_pp_it_7 ) : ( n252 ) ;
assign n254 =  ( n4 ) ? ( gb_pp_it_8 ) : ( n253 ) ;
assign n255 =  ( n28 ) ? ( gb_pp_it_9 ) : ( gb_pp_it_9 ) ;
assign n256 =  ( n25 ) ? ( gb_pp_it_9 ) : ( n255 ) ;
assign n257 =  ( n20 ) ? ( gb_pp_it_9 ) : ( n256 ) ;
assign n258 =  ( n13 ) ? ( gb_pp_it_8 ) : ( n257 ) ;
assign n259 =  ( n4 ) ? ( gb_pp_it_9 ) : ( n258 ) ;
assign n260 =  ( n28 ) ? ( LB1D_uIn ) : ( in_stream_buff_0 ) ;
assign n261 =  ( n25 ) ? ( in_stream_buff_0 ) : ( n260 ) ;
assign n262 =  ( n20 ) ? ( in_stream_buff_0 ) : ( n261 ) ;
assign n263 =  ( n13 ) ? ( in_stream_buff_0 ) : ( n262 ) ;
assign n264 =  ( n4 ) ? ( in_stream_buff_0 ) : ( n263 ) ;
assign n265 =  ( n28 ) ? ( in_stream_buff_0 ) : ( in_stream_buff_1 ) ;
assign n266 =  ( n25 ) ? ( in_stream_buff_1 ) : ( n265 ) ;
assign n267 =  ( n20 ) ? ( in_stream_buff_1 ) : ( n266 ) ;
assign n268 =  ( n13 ) ? ( in_stream_buff_1 ) : ( n267 ) ;
assign n269 =  ( n4 ) ? ( in_stream_buff_1 ) : ( n268 ) ;
assign n270 =  ( in_stream_full ) == ( 1'd1 )  ;
assign n271 =  ( n270 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n272 =  ( n28 ) ? ( 1'd0 ) : ( in_stream_empty ) ;
assign n273 =  ( n25 ) ? ( n271 ) : ( n272 ) ;
assign n274 =  ( n20 ) ? ( in_stream_empty ) : ( n273 ) ;
assign n275 =  ( n13 ) ? ( in_stream_empty ) : ( n274 ) ;
assign n276 =  ( n4 ) ? ( in_stream_empty ) : ( n275 ) ;
assign n277 =  ( in_stream_empty ) == ( 1'd1 )  ;
assign n278 =  ( n277 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n279 =  ( n28 ) ? ( n278 ) : ( in_stream_full ) ;
assign n280 =  ( n25 ) ? ( 1'd0 ) : ( n279 ) ;
assign n281 =  ( n20 ) ? ( in_stream_full ) : ( n280 ) ;
assign n282 =  ( n13 ) ? ( in_stream_full ) : ( n281 ) ;
assign n283 =  ( n4 ) ? ( in_stream_full ) : ( n282 ) ;
assign n284 =  ( n270 ) ? ( in_stream_buff_1 ) : ( in_stream_buff_0 ) ;
assign n285 =  ( LB2D_proc_w ) == ( 64'd0 )  ;
assign n286 =  ( LB2D_proc_x ) - ( 9'd1 )  ;
assign n287 =  (  LB2D_proc_7 [ n286 ] )  ;
assign n288 =  ( LB2D_proc_w ) == ( 64'd1 )  ;
assign n289 =  (  LB2D_proc_0 [ n286 ] )  ;
assign n290 =  ( LB2D_proc_w ) == ( 64'd2 )  ;
assign n291 =  (  LB2D_proc_1 [ n286 ] )  ;
assign n292 =  ( LB2D_proc_w ) == ( 64'd3 )  ;
assign n293 =  (  LB2D_proc_2 [ n286 ] )  ;
assign n294 =  ( LB2D_proc_w ) == ( 64'd4 )  ;
assign n295 =  (  LB2D_proc_3 [ n286 ] )  ;
assign n296 =  ( LB2D_proc_w ) == ( 64'd5 )  ;
assign n297 =  (  LB2D_proc_4 [ n286 ] )  ;
assign n298 =  ( LB2D_proc_w ) == ( 64'd6 )  ;
assign n299 =  (  LB2D_proc_5 [ n286 ] )  ;
assign n300 =  (  LB2D_proc_6 [ n286 ] )  ;
assign n301 =  ( n298 ) ? ( n299 ) : ( n300 ) ;
assign n302 =  ( n296 ) ? ( n297 ) : ( n301 ) ;
assign n303 =  ( n294 ) ? ( n295 ) : ( n302 ) ;
assign n304 =  ( n292 ) ? ( n293 ) : ( n303 ) ;
assign n305 =  ( n290 ) ? ( n291 ) : ( n304 ) ;
assign n306 =  ( n288 ) ? ( n289 ) : ( n305 ) ;
assign n307 =  ( n285 ) ? ( n287 ) : ( n306 ) ;
assign n308 =  ( n298 ) ? ( n297 ) : ( n299 ) ;
assign n309 =  ( n296 ) ? ( n295 ) : ( n308 ) ;
assign n310 =  ( n294 ) ? ( n293 ) : ( n309 ) ;
assign n311 =  ( n292 ) ? ( n291 ) : ( n310 ) ;
assign n312 =  ( n290 ) ? ( n289 ) : ( n311 ) ;
assign n313 =  ( n288 ) ? ( n287 ) : ( n312 ) ;
assign n314 =  ( n285 ) ? ( n300 ) : ( n313 ) ;
assign n315 =  ( n298 ) ? ( n295 ) : ( n297 ) ;
assign n316 =  ( n296 ) ? ( n293 ) : ( n315 ) ;
assign n317 =  ( n294 ) ? ( n291 ) : ( n316 ) ;
assign n318 =  ( n292 ) ? ( n289 ) : ( n317 ) ;
assign n319 =  ( n290 ) ? ( n287 ) : ( n318 ) ;
assign n320 =  ( n288 ) ? ( n300 ) : ( n319 ) ;
assign n321 =  ( n285 ) ? ( n299 ) : ( n320 ) ;
assign n322 =  ( n298 ) ? ( n293 ) : ( n295 ) ;
assign n323 =  ( n296 ) ? ( n291 ) : ( n322 ) ;
assign n324 =  ( n294 ) ? ( n289 ) : ( n323 ) ;
assign n325 =  ( n292 ) ? ( n287 ) : ( n324 ) ;
assign n326 =  ( n290 ) ? ( n300 ) : ( n325 ) ;
assign n327 =  ( n288 ) ? ( n299 ) : ( n326 ) ;
assign n328 =  ( n285 ) ? ( n297 ) : ( n327 ) ;
assign n329 =  ( n298 ) ? ( n291 ) : ( n293 ) ;
assign n330 =  ( n296 ) ? ( n289 ) : ( n329 ) ;
assign n331 =  ( n294 ) ? ( n287 ) : ( n330 ) ;
assign n332 =  ( n292 ) ? ( n300 ) : ( n331 ) ;
assign n333 =  ( n290 ) ? ( n299 ) : ( n332 ) ;
assign n334 =  ( n288 ) ? ( n297 ) : ( n333 ) ;
assign n335 =  ( n285 ) ? ( n295 ) : ( n334 ) ;
assign n336 =  ( n298 ) ? ( n289 ) : ( n291 ) ;
assign n337 =  ( n296 ) ? ( n287 ) : ( n336 ) ;
assign n338 =  ( n294 ) ? ( n300 ) : ( n337 ) ;
assign n339 =  ( n292 ) ? ( n299 ) : ( n338 ) ;
assign n340 =  ( n290 ) ? ( n297 ) : ( n339 ) ;
assign n341 =  ( n288 ) ? ( n295 ) : ( n340 ) ;
assign n342 =  ( n285 ) ? ( n293 ) : ( n341 ) ;
assign n343 =  ( n298 ) ? ( n287 ) : ( n289 ) ;
assign n344 =  ( n296 ) ? ( n300 ) : ( n343 ) ;
assign n345 =  ( n294 ) ? ( n299 ) : ( n344 ) ;
assign n346 =  ( n292 ) ? ( n297 ) : ( n345 ) ;
assign n347 =  ( n290 ) ? ( n295 ) : ( n346 ) ;
assign n348 =  ( n288 ) ? ( n293 ) : ( n347 ) ;
assign n349 =  ( n285 ) ? ( n291 ) : ( n348 ) ;
assign n350 =  ( n298 ) ? ( n300 ) : ( n287 ) ;
assign n351 =  ( n296 ) ? ( n299 ) : ( n350 ) ;
assign n352 =  ( n294 ) ? ( n297 ) : ( n351 ) ;
assign n353 =  ( n292 ) ? ( n295 ) : ( n352 ) ;
assign n354 =  ( n290 ) ? ( n293 ) : ( n353 ) ;
assign n355 =  ( n288 ) ? ( n291 ) : ( n354 ) ;
assign n356 =  ( n285 ) ? ( n289 ) : ( n355 ) ;
assign n357 =  { ( n349 ) , ( n356 ) }  ;
assign n358 =  { ( n342 ) , ( n357 ) }  ;
assign n359 =  { ( n335 ) , ( n358 ) }  ;
assign n360 =  { ( n328 ) , ( n359 ) }  ;
assign n361 =  { ( n321 ) , ( n360 ) }  ;
assign n362 =  { ( n314 ) , ( n361 ) }  ;
assign n363 =  { ( n307 ) , ( n362 ) }  ;
assign n364 =  { ( n284 ) , ( n363 ) }  ;
assign n365 =  ( n23 ) ? ( slice_stream_buff_0 ) : ( n364 ) ;
assign n366 =  ( n28 ) ? ( slice_stream_buff_0 ) : ( slice_stream_buff_0 ) ;
assign n367 =  ( n25 ) ? ( n365 ) : ( n366 ) ;
assign n368 =  ( n20 ) ? ( slice_stream_buff_0 ) : ( n367 ) ;
assign n369 =  ( n13 ) ? ( slice_stream_buff_0 ) : ( n368 ) ;
assign n370 =  ( n4 ) ? ( slice_stream_buff_0 ) : ( n369 ) ;
assign n371 =  ( n23 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n372 =  ( n28 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_1 ) ;
assign n373 =  ( n25 ) ? ( n371 ) : ( n372 ) ;
assign n374 =  ( n20 ) ? ( slice_stream_buff_1 ) : ( n373 ) ;
assign n375 =  ( n13 ) ? ( slice_stream_buff_1 ) : ( n374 ) ;
assign n376 =  ( n4 ) ? ( slice_stream_buff_1 ) : ( n375 ) ;
assign n377 =  ( n116 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n378 =  ( n23 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n379 =  ( n28 ) ? ( slice_stream_empty ) : ( slice_stream_empty ) ;
assign n380 =  ( n25 ) ? ( n378 ) : ( n379 ) ;
assign n381 =  ( n20 ) ? ( n377 ) : ( n380 ) ;
assign n382 =  ( n13 ) ? ( slice_stream_empty ) : ( n381 ) ;
assign n383 =  ( n4 ) ? ( slice_stream_empty ) : ( n382 ) ;
assign n384 =  ( slice_stream_empty ) == ( 1'd1 )  ;
assign n385 =  ( n384 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n386 =  ( n23 ) ? ( 1'd0 ) : ( n385 ) ;
assign n387 =  ( n28 ) ? ( slice_stream_full ) : ( slice_stream_full ) ;
assign n388 =  ( n25 ) ? ( n386 ) : ( n387 ) ;
assign n389 =  ( n20 ) ? ( 1'd0 ) : ( n388 ) ;
assign n390 =  ( n13 ) ? ( slice_stream_full ) : ( n389 ) ;
assign n391 =  ( n4 ) ? ( slice_stream_full ) : ( n390 ) ;
assign n392 =  ( LB2D_shift_x ) >= ( 9'd8 )  ;
assign n393 =  ( LB2D_shift_x ) == ( 9'd0 )  ;
assign n394 =  ( n392 ) | ( n393 )  ;
assign n395 = n117[71:64] ;
assign n396 = LB2D_shift_7[71:64] ;
assign n397 = LB2D_shift_6[71:64] ;
assign n398 = LB2D_shift_5[71:64] ;
assign n399 = LB2D_shift_4[71:64] ;
assign n400 = LB2D_shift_3[71:64] ;
assign n401 = LB2D_shift_2[71:64] ;
assign n402 = LB2D_shift_1[71:64] ;
assign n403 = LB2D_shift_0[71:64] ;
assign n404 =  { ( n402 ) , ( n403 ) }  ;
assign n405 =  { ( n401 ) , ( n404 ) }  ;
assign n406 =  { ( n400 ) , ( n405 ) }  ;
assign n407 =  { ( n399 ) , ( n406 ) }  ;
assign n408 =  { ( n398 ) , ( n407 ) }  ;
assign n409 =  { ( n397 ) , ( n408 ) }  ;
assign n410 =  { ( n396 ) , ( n409 ) }  ;
assign n411 =  { ( n395 ) , ( n410 ) }  ;
assign n412 = n117[63:56] ;
assign n413 = LB2D_shift_7[63:56] ;
assign n414 = LB2D_shift_6[63:56] ;
assign n415 = LB2D_shift_5[63:56] ;
assign n416 = LB2D_shift_4[63:56] ;
assign n417 = LB2D_shift_3[63:56] ;
assign n418 = LB2D_shift_2[63:56] ;
assign n419 = LB2D_shift_1[63:56] ;
assign n420 = LB2D_shift_0[63:56] ;
assign n421 =  { ( n419 ) , ( n420 ) }  ;
assign n422 =  { ( n418 ) , ( n421 ) }  ;
assign n423 =  { ( n417 ) , ( n422 ) }  ;
assign n424 =  { ( n416 ) , ( n423 ) }  ;
assign n425 =  { ( n415 ) , ( n424 ) }  ;
assign n426 =  { ( n414 ) , ( n425 ) }  ;
assign n427 =  { ( n413 ) , ( n426 ) }  ;
assign n428 =  { ( n412 ) , ( n427 ) }  ;
assign n429 = n117[55:48] ;
assign n430 = LB2D_shift_7[55:48] ;
assign n431 = LB2D_shift_6[55:48] ;
assign n432 = LB2D_shift_5[55:48] ;
assign n433 = LB2D_shift_4[55:48] ;
assign n434 = LB2D_shift_3[55:48] ;
assign n435 = LB2D_shift_2[55:48] ;
assign n436 = LB2D_shift_1[55:48] ;
assign n437 = LB2D_shift_0[55:48] ;
assign n438 =  { ( n436 ) , ( n437 ) }  ;
assign n439 =  { ( n435 ) , ( n438 ) }  ;
assign n440 =  { ( n434 ) , ( n439 ) }  ;
assign n441 =  { ( n433 ) , ( n440 ) }  ;
assign n442 =  { ( n432 ) , ( n441 ) }  ;
assign n443 =  { ( n431 ) , ( n442 ) }  ;
assign n444 =  { ( n430 ) , ( n443 ) }  ;
assign n445 =  { ( n429 ) , ( n444 ) }  ;
assign n446 = n117[47:40] ;
assign n447 = LB2D_shift_7[47:40] ;
assign n448 = LB2D_shift_6[47:40] ;
assign n449 = LB2D_shift_5[47:40] ;
assign n450 = LB2D_shift_4[47:40] ;
assign n451 = LB2D_shift_3[47:40] ;
assign n452 = LB2D_shift_2[47:40] ;
assign n453 = LB2D_shift_1[47:40] ;
assign n454 = LB2D_shift_0[47:40] ;
assign n455 =  { ( n453 ) , ( n454 ) }  ;
assign n456 =  { ( n452 ) , ( n455 ) }  ;
assign n457 =  { ( n451 ) , ( n456 ) }  ;
assign n458 =  { ( n450 ) , ( n457 ) }  ;
assign n459 =  { ( n449 ) , ( n458 ) }  ;
assign n460 =  { ( n448 ) , ( n459 ) }  ;
assign n461 =  { ( n447 ) , ( n460 ) }  ;
assign n462 =  { ( n446 ) , ( n461 ) }  ;
assign n463 = n117[39:32] ;
assign n464 = LB2D_shift_7[39:32] ;
assign n465 = LB2D_shift_6[39:32] ;
assign n466 = LB2D_shift_5[39:32] ;
assign n467 = LB2D_shift_4[39:32] ;
assign n468 = LB2D_shift_3[39:32] ;
assign n469 = LB2D_shift_2[39:32] ;
assign n470 = LB2D_shift_1[39:32] ;
assign n471 = LB2D_shift_0[39:32] ;
assign n472 =  { ( n470 ) , ( n471 ) }  ;
assign n473 =  { ( n469 ) , ( n472 ) }  ;
assign n474 =  { ( n468 ) , ( n473 ) }  ;
assign n475 =  { ( n467 ) , ( n474 ) }  ;
assign n476 =  { ( n466 ) , ( n475 ) }  ;
assign n477 =  { ( n465 ) , ( n476 ) }  ;
assign n478 =  { ( n464 ) , ( n477 ) }  ;
assign n479 =  { ( n463 ) , ( n478 ) }  ;
assign n480 = n117[31:24] ;
assign n481 = LB2D_shift_7[31:24] ;
assign n482 = LB2D_shift_6[31:24] ;
assign n483 = LB2D_shift_5[31:24] ;
assign n484 = LB2D_shift_4[31:24] ;
assign n485 = LB2D_shift_3[31:24] ;
assign n486 = LB2D_shift_2[31:24] ;
assign n487 = LB2D_shift_1[31:24] ;
assign n488 = LB2D_shift_0[31:24] ;
assign n489 =  { ( n487 ) , ( n488 ) }  ;
assign n490 =  { ( n486 ) , ( n489 ) }  ;
assign n491 =  { ( n485 ) , ( n490 ) }  ;
assign n492 =  { ( n484 ) , ( n491 ) }  ;
assign n493 =  { ( n483 ) , ( n492 ) }  ;
assign n494 =  { ( n482 ) , ( n493 ) }  ;
assign n495 =  { ( n481 ) , ( n494 ) }  ;
assign n496 =  { ( n480 ) , ( n495 ) }  ;
assign n497 = n117[23:16] ;
assign n498 = LB2D_shift_7[23:16] ;
assign n499 = LB2D_shift_6[23:16] ;
assign n500 = LB2D_shift_5[23:16] ;
assign n501 = LB2D_shift_4[23:16] ;
assign n502 = LB2D_shift_3[23:16] ;
assign n503 = LB2D_shift_2[23:16] ;
assign n504 = LB2D_shift_1[23:16] ;
assign n505 = LB2D_shift_0[23:16] ;
assign n506 =  { ( n504 ) , ( n505 ) }  ;
assign n507 =  { ( n503 ) , ( n506 ) }  ;
assign n508 =  { ( n502 ) , ( n507 ) }  ;
assign n509 =  { ( n501 ) , ( n508 ) }  ;
assign n510 =  { ( n500 ) , ( n509 ) }  ;
assign n511 =  { ( n499 ) , ( n510 ) }  ;
assign n512 =  { ( n498 ) , ( n511 ) }  ;
assign n513 =  { ( n497 ) , ( n512 ) }  ;
assign n514 = n117[15:8] ;
assign n515 = LB2D_shift_7[15:8] ;
assign n516 = LB2D_shift_6[15:8] ;
assign n517 = LB2D_shift_5[15:8] ;
assign n518 = LB2D_shift_4[15:8] ;
assign n519 = LB2D_shift_3[15:8] ;
assign n520 = LB2D_shift_2[15:8] ;
assign n521 = LB2D_shift_1[15:8] ;
assign n522 = LB2D_shift_0[15:8] ;
assign n523 =  { ( n521 ) , ( n522 ) }  ;
assign n524 =  { ( n520 ) , ( n523 ) }  ;
assign n525 =  { ( n519 ) , ( n524 ) }  ;
assign n526 =  { ( n518 ) , ( n525 ) }  ;
assign n527 =  { ( n517 ) , ( n526 ) }  ;
assign n528 =  { ( n516 ) , ( n527 ) }  ;
assign n529 =  { ( n515 ) , ( n528 ) }  ;
assign n530 =  { ( n514 ) , ( n529 ) }  ;
assign n531 = n117[7:0] ;
assign n532 = LB2D_shift_7[7:0] ;
assign n533 = LB2D_shift_6[7:0] ;
assign n534 = LB2D_shift_5[7:0] ;
assign n535 = LB2D_shift_4[7:0] ;
assign n536 = LB2D_shift_3[7:0] ;
assign n537 = LB2D_shift_2[7:0] ;
assign n538 = LB2D_shift_1[7:0] ;
assign n539 = LB2D_shift_0[7:0] ;
assign n540 =  { ( n538 ) , ( n539 ) }  ;
assign n541 =  { ( n537 ) , ( n540 ) }  ;
assign n542 =  { ( n536 ) , ( n541 ) }  ;
assign n543 =  { ( n535 ) , ( n542 ) }  ;
assign n544 =  { ( n534 ) , ( n543 ) }  ;
assign n545 =  { ( n533 ) , ( n544 ) }  ;
assign n546 =  { ( n532 ) , ( n545 ) }  ;
assign n547 =  { ( n531 ) , ( n546 ) }  ;
assign n548 =  { ( n530 ) , ( n547 ) }  ;
assign n549 =  { ( n513 ) , ( n548 ) }  ;
assign n550 =  { ( n496 ) , ( n549 ) }  ;
assign n551 =  { ( n479 ) , ( n550 ) }  ;
assign n552 =  { ( n462 ) , ( n551 ) }  ;
assign n553 =  { ( n445 ) , ( n552 ) }  ;
assign n554 =  { ( n428 ) , ( n553 ) }  ;
assign n555 =  { ( n411 ) , ( n554 ) }  ;
assign n556 =  ( n394 ) ? ( n555 ) : ( stencil_stream_buff_0 ) ;
assign n557 =  ( n28 ) ? ( stencil_stream_buff_0 ) : ( stencil_stream_buff_0 ) ;
assign n558 =  ( n25 ) ? ( stencil_stream_buff_0 ) : ( n557 ) ;
assign n559 =  ( n20 ) ? ( n556 ) : ( n558 ) ;
assign n560 =  ( n13 ) ? ( stencil_stream_buff_0 ) : ( n559 ) ;
assign n561 =  ( n4 ) ? ( stencil_stream_buff_0 ) : ( n560 ) ;
assign n562 =  ( n20 ) & ( n394 )  ;
assign n563 =  ( n28 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_1 ) ;
assign n564 =  ( n25 ) ? ( stencil_stream_buff_1 ) : ( n563 ) ;
assign n565 =  ( n562 ) ? ( stencil_stream_buff_0 ) : ( n564 ) ;
assign n566 =  ( n13 ) ? ( stencil_stream_buff_1 ) : ( n565 ) ;
assign n567 =  ( n4 ) ? ( stencil_stream_buff_1 ) : ( n566 ) ;
assign n568 =  ( n141 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n569 = ~ ( n394 ) ;
assign n570 =  ( n569 ) ? ( stencil_stream_empty ) : ( 1'd0 ) ;
assign n571 =  ( n28 ) ? ( stencil_stream_empty ) : ( stencil_stream_empty ) ;
assign n572 =  ( n25 ) ? ( stencil_stream_empty ) : ( n571 ) ;
assign n573 =  ( n20 ) ? ( n570 ) : ( n572 ) ;
assign n574 =  ( n13 ) ? ( n568 ) : ( n573 ) ;
assign n575 =  ( n4 ) ? ( stencil_stream_empty ) : ( n574 ) ;
assign n576 =  ( n9 ) ? ( 1'd0 ) : ( 1'd0 ) ;
assign n577 =  ( stencil_stream_empty ) == ( 1'd1 )  ;
assign n578 =  ( n577 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n579 =  ( n569 ) ? ( stencil_stream_full ) : ( n578 ) ;
assign n580 =  ( n28 ) ? ( stencil_stream_full ) : ( stencil_stream_full ) ;
assign n581 =  ( n25 ) ? ( stencil_stream_full ) : ( n580 ) ;
assign n582 =  ( n20 ) ? ( n579 ) : ( n581 ) ;
assign n583 =  ( n13 ) ? ( n576 ) : ( n582 ) ;
assign n584 =  ( n4 ) ? ( stencil_stream_full ) : ( n583 ) ;
assign n585 = ~ ( n4 ) ;
assign n586 =  ( 1'b1 ) & ( n585 )  ;
assign n587 = ~ ( n13 ) ;
assign n588 =  ( n586 ) & ( n587 )  ;
assign n589 = ~ ( n20 ) ;
assign n590 =  ( n588 ) & ( n589 )  ;
assign n591 = ~ ( n25 ) ;
assign n592 =  ( n590 ) & ( n591 )  ;
assign n593 = ~ ( n28 ) ;
assign n594 =  ( n592 ) & ( n593 )  ;
assign n595 =  ( n592 ) & ( n28 )  ;
assign n596 =  ( n590 ) & ( n25 )  ;
assign n597 = ~ ( n285 ) ;
assign n598 =  ( n596 ) & ( n597 )  ;
assign n599 =  ( n596 ) & ( n285 )  ;
assign n600 =  ( n588 ) & ( n20 )  ;
assign n601 =  ( n586 ) & ( n13 )  ;
assign n602 =  ( 1'b1 ) & ( n4 )  ;
assign LB2D_proc_0_addr0 = n599 ? (n286) : (0);
assign LB2D_proc_0_data0 = n599 ? (n284) : ('dx);
assign LB2D_proc_0_wen0 = n599 ? ( 1'b1 ) : (1'b0);
assign n603 = ~ ( n288 ) ;
assign n604 =  ( n596 ) & ( n603 )  ;
assign n605 =  ( n596 ) & ( n288 )  ;
assign LB2D_proc_1_addr0 = n605 ? (n286) : (0);
assign LB2D_proc_1_data0 = n605 ? (n284) : ('dx);
assign LB2D_proc_1_wen0 = n605 ? ( 1'b1 ) : (1'b0);
assign n606 = ~ ( n290 ) ;
assign n607 =  ( n596 ) & ( n606 )  ;
assign n608 =  ( n596 ) & ( n290 )  ;
assign LB2D_proc_2_addr0 = n608 ? (n286) : (0);
assign LB2D_proc_2_data0 = n608 ? (n284) : ('dx);
assign LB2D_proc_2_wen0 = n608 ? ( 1'b1 ) : (1'b0);
assign n609 = ~ ( n292 ) ;
assign n610 =  ( n596 ) & ( n609 )  ;
assign n611 =  ( n596 ) & ( n292 )  ;
assign LB2D_proc_3_addr0 = n611 ? (n286) : (0);
assign LB2D_proc_3_data0 = n611 ? (n284) : ('dx);
assign LB2D_proc_3_wen0 = n611 ? ( 1'b1 ) : (1'b0);
assign n612 = ~ ( n294 ) ;
assign n613 =  ( n596 ) & ( n612 )  ;
assign n614 =  ( n596 ) & ( n294 )  ;
assign LB2D_proc_4_addr0 = n614 ? (n286) : (0);
assign LB2D_proc_4_data0 = n614 ? (n284) : ('dx);
assign LB2D_proc_4_wen0 = n614 ? ( 1'b1 ) : (1'b0);
assign n615 = ~ ( n296 ) ;
assign n616 =  ( n596 ) & ( n615 )  ;
assign n617 =  ( n596 ) & ( n296 )  ;
assign LB2D_proc_5_addr0 = n617 ? (n286) : (0);
assign LB2D_proc_5_data0 = n617 ? (n284) : ('dx);
assign LB2D_proc_5_wen0 = n617 ? ( 1'b1 ) : (1'b0);
assign n618 = ~ ( n298 ) ;
assign n619 =  ( n596 ) & ( n618 )  ;
assign n620 =  ( n596 ) & ( n298 )  ;
assign LB2D_proc_6_addr0 = n620 ? (n286) : (0);
assign LB2D_proc_6_data0 = n620 ? (n284) : ('dx);
assign LB2D_proc_6_wen0 = n620 ? ( 1'b1 ) : (1'b0);
assign n621 = ~ ( n56 ) ;
assign n622 =  ( n596 ) & ( n621 )  ;
assign n623 =  ( n596 ) & ( n56 )  ;
assign LB2D_proc_7_addr0 = n623 ? (n286) : (0);
assign LB2D_proc_7_data0 = n623 ? (n284) : ('dx);
assign LB2D_proc_7_wen0 = n623 ? ( 1'b1 ) : (1'b0);
always @(posedge clk) begin
   if(rst) begin
       LB1D_buff <= LB1D_buff;
       LB1D_in <= LB1D_in;
       LB1D_it_1 <= LB1D_it_1;
       LB1D_p_cnt <= LB1D_p_cnt;
       LB1D_uIn <= LB1D_uIn;
       LB2D_proc_w <= LB2D_proc_w;
       LB2D_proc_x <= LB2D_proc_x;
       LB2D_proc_y <= LB2D_proc_y;
       LB2D_shift_0 <= LB2D_shift_0;
       LB2D_shift_1 <= LB2D_shift_1;
       LB2D_shift_2 <= LB2D_shift_2;
       LB2D_shift_3 <= LB2D_shift_3;
       LB2D_shift_4 <= LB2D_shift_4;
       LB2D_shift_5 <= LB2D_shift_5;
       LB2D_shift_6 <= LB2D_shift_6;
       LB2D_shift_7 <= LB2D_shift_7;
       LB2D_shift_x <= LB2D_shift_x;
       LB2D_shift_y <= LB2D_shift_y;
       arg_0_TDATA <= arg_0_TDATA;
       arg_0_TVALID <= arg_0_TVALID;
       arg_1_TREADY <= arg_1_TREADY;
       gb_exit_it_1 <= gb_exit_it_1;
       gb_exit_it_2 <= gb_exit_it_2;
       gb_exit_it_3 <= gb_exit_it_3;
       gb_exit_it_4 <= gb_exit_it_4;
       gb_exit_it_5 <= gb_exit_it_5;
       gb_exit_it_6 <= gb_exit_it_6;
       gb_exit_it_7 <= gb_exit_it_7;
       gb_exit_it_8 <= gb_exit_it_8;
       gb_p_cnt <= gb_p_cnt;
       gb_pp_it_1 <= gb_pp_it_1;
       gb_pp_it_2 <= gb_pp_it_2;
       gb_pp_it_3 <= gb_pp_it_3;
       gb_pp_it_4 <= gb_pp_it_4;
       gb_pp_it_5 <= gb_pp_it_5;
       gb_pp_it_6 <= gb_pp_it_6;
       gb_pp_it_7 <= gb_pp_it_7;
       gb_pp_it_8 <= gb_pp_it_8;
       gb_pp_it_9 <= gb_pp_it_9;
       in_stream_buff_0 <= in_stream_buff_0;
       in_stream_buff_1 <= in_stream_buff_1;
       in_stream_empty <= in_stream_empty;
       in_stream_full <= in_stream_full;
       slice_stream_buff_0 <= slice_stream_buff_0;
       slice_stream_buff_1 <= slice_stream_buff_1;
       slice_stream_empty <= slice_stream_empty;
       slice_stream_full <= slice_stream_full;
       stencil_stream_buff_0 <= stencil_stream_buff_0;
       stencil_stream_buff_1 <= stencil_stream_buff_1;
       stencil_stream_empty <= stencil_stream_empty;
       stencil_stream_full <= stencil_stream_full;
   end
   else if(step) begin
       LB1D_buff <= n33;
       LB1D_in <= n38;
       LB1D_it_1 <= n43;
       LB1D_p_cnt <= n50;
       LB1D_uIn <= n54;
       LB2D_proc_w <= n64;
       LB2D_proc_x <= n71;
       LB2D_proc_y <= n80;
       LB2D_shift_0 <= n85;
       LB2D_shift_1 <= n90;
       LB2D_shift_2 <= n95;
       LB2D_shift_3 <= n100;
       LB2D_shift_4 <= n105;
       LB2D_shift_5 <= n110;
       LB2D_shift_6 <= n115;
       LB2D_shift_7 <= n122;
       LB2D_shift_x <= n130;
       LB2D_shift_y <= n140;
       arg_0_TDATA <= n150;
       arg_0_TVALID <= n159;
       arg_1_TREADY <= n164;
       gb_exit_it_1 <= n171;
       gb_exit_it_2 <= n176;
       gb_exit_it_3 <= n181;
       gb_exit_it_4 <= n186;
       gb_exit_it_5 <= n191;
       gb_exit_it_6 <= n196;
       gb_exit_it_7 <= n201;
       gb_exit_it_8 <= n206;
       gb_p_cnt <= n214;
       gb_pp_it_1 <= n219;
       gb_pp_it_2 <= n224;
       gb_pp_it_3 <= n229;
       gb_pp_it_4 <= n234;
       gb_pp_it_5 <= n239;
       gb_pp_it_6 <= n244;
       gb_pp_it_7 <= n249;
       gb_pp_it_8 <= n254;
       gb_pp_it_9 <= n259;
       in_stream_buff_0 <= n264;
       in_stream_buff_1 <= n269;
       in_stream_empty <= n276;
       in_stream_full <= n283;
       slice_stream_buff_0 <= n370;
       slice_stream_buff_1 <= n376;
       slice_stream_empty <= n383;
       slice_stream_full <= n391;
       stencil_stream_buff_0 <= n561;
       stencil_stream_buff_1 <= n567;
       stencil_stream_empty <= n575;
       stencil_stream_full <= n584;
       if (LB2D_proc_0_wen0) begin
           LB2D_proc_0 [ LB2D_proc_0_addr0 ] <= LB2D_proc_0_data0 ;
       end
       if (LB2D_proc_1_wen0) begin
           LB2D_proc_1 [ LB2D_proc_1_addr0 ] <= LB2D_proc_1_data0 ;
       end
       if (LB2D_proc_2_wen0) begin
           LB2D_proc_2 [ LB2D_proc_2_addr0 ] <= LB2D_proc_2_data0 ;
       end
       if (LB2D_proc_3_wen0) begin
           LB2D_proc_3 [ LB2D_proc_3_addr0 ] <= LB2D_proc_3_data0 ;
       end
       if (LB2D_proc_4_wen0) begin
           LB2D_proc_4 [ LB2D_proc_4_addr0 ] <= LB2D_proc_4_data0 ;
       end
       if (LB2D_proc_5_wen0) begin
           LB2D_proc_5 [ LB2D_proc_5_addr0 ] <= LB2D_proc_5_data0 ;
       end
       if (LB2D_proc_6_wen0) begin
           LB2D_proc_6 [ LB2D_proc_6_addr0 ] <= LB2D_proc_6_data0 ;
       end
       if (LB2D_proc_7_wen0) begin
           LB2D_proc_7 [ LB2D_proc_7_addr0 ] <= LB2D_proc_7_data0 ;
       end
   end
end
endmodule
