module GB(
arg_0_TREADY,
arg_1_TDATA,
arg_1_TVALID,
LB1D_buff,
LB1D_in,
LB1D_it_1,
LB1D_p_cnt,
LB2D_proc_w,
LB2D_proc_x,
LB2D_proc_y,
LB2D_shift_0,
LB2D_shift_1,
LB2D_shift_2,
LB2D_shift_3,
LB2D_shift_4,
LB2D_shift_5,
LB2D_shift_6,
LB2D_shift_7,
LB2D_shift_x,
LB2D_shift_y,
arg_0_TDATA,
arg_0_TVALID,
arg_1_TREADY,
gb_exit_it_1,
gb_exit_it_2,
gb_exit_it_3,
gb_exit_it_4,
gb_exit_it_5,
gb_exit_it_6,
gb_exit_it_7,
gb_exit_it_8,
gb_p_cnt,
gb_pp_it_1,
gb_pp_it_2,
gb_pp_it_3,
gb_pp_it_4,
gb_pp_it_5,
gb_pp_it_6,
gb_pp_it_7,
gb_pp_it_8,
gb_pp_it_9,
in_stream_buff_0,
in_stream_buff_1,
in_stream_empty,
in_stream_full,
slice_stream_buff_0,
slice_stream_buff_1,
slice_stream_empty,
slice_stream_full,
stencil_stream_buff_0,
stencil_stream_buff_1,
stencil_stream_empty,
stencil_stream_full,
clk,rst,
step
);
input            arg_0_TREADY;
input      [7:0] arg_1_TDATA;
input            arg_1_TVALID;
input clk;
input rst;
input step;
output      [7:0] LB1D_buff;
output      [7:0] LB1D_in;
output            LB1D_it_1;
output     [18:0] LB1D_p_cnt;
output     [63:0] LB2D_proc_w;
output      [8:0] LB2D_proc_x;
output      [9:0] LB2D_proc_y;
output     [71:0] LB2D_shift_0;
output     [71:0] LB2D_shift_1;
output     [71:0] LB2D_shift_2;
output     [71:0] LB2D_shift_3;
output     [71:0] LB2D_shift_4;
output     [71:0] LB2D_shift_5;
output     [71:0] LB2D_shift_6;
output     [71:0] LB2D_shift_7;
output      [8:0] LB2D_shift_x;
output      [9:0] LB2D_shift_y;
output      [7:0] arg_0_TDATA;
output            arg_0_TVALID;
output            arg_1_TREADY;
output            gb_exit_it_1;
output            gb_exit_it_2;
output            gb_exit_it_3;
output            gb_exit_it_4;
output            gb_exit_it_5;
output            gb_exit_it_6;
output            gb_exit_it_7;
output            gb_exit_it_8;
output     [18:0] gb_p_cnt;
output            gb_pp_it_1;
output            gb_pp_it_2;
output            gb_pp_it_3;
output            gb_pp_it_4;
output            gb_pp_it_5;
output            gb_pp_it_6;
output            gb_pp_it_7;
output            gb_pp_it_8;
output            gb_pp_it_9;
output      [7:0] in_stream_buff_0;
output      [7:0] in_stream_buff_1;
output            in_stream_empty;
output            in_stream_full;
output     [71:0] slice_stream_buff_0;
output     [71:0] slice_stream_buff_1;
output            slice_stream_empty;
output            slice_stream_full;
output    [647:0] stencil_stream_buff_0;
output    [647:0] stencil_stream_buff_1;
output            stencil_stream_empty;
output            stencil_stream_full;
reg      [7:0] LB1D_buff;
reg      [7:0] LB1D_in;
reg            LB1D_it_1;
reg     [18:0] LB1D_p_cnt;
reg     [63:0] LB2D_proc_w;
reg      [8:0] LB2D_proc_x;
reg      [9:0] LB2D_proc_y;
reg     [71:0] LB2D_shift_0;
reg     [71:0] LB2D_shift_1;
reg     [71:0] LB2D_shift_2;
reg     [71:0] LB2D_shift_3;
reg     [71:0] LB2D_shift_4;
reg     [71:0] LB2D_shift_5;
reg     [71:0] LB2D_shift_6;
reg     [71:0] LB2D_shift_7;
reg      [8:0] LB2D_shift_x;
reg      [9:0] LB2D_shift_y;
reg      [7:0] arg_0_TDATA;
reg            arg_0_TVALID;
reg            arg_1_TREADY;
reg            gb_exit_it_1;
reg            gb_exit_it_2;
reg            gb_exit_it_3;
reg            gb_exit_it_4;
reg            gb_exit_it_5;
reg            gb_exit_it_6;
reg            gb_exit_it_7;
reg            gb_exit_it_8;
reg     [18:0] gb_p_cnt;
reg            gb_pp_it_1;
reg            gb_pp_it_2;
reg            gb_pp_it_3;
reg            gb_pp_it_4;
reg            gb_pp_it_5;
reg            gb_pp_it_6;
reg            gb_pp_it_7;
reg            gb_pp_it_8;
reg            gb_pp_it_9;
reg      [7:0] in_stream_buff_0;
reg      [7:0] in_stream_buff_1;
reg            in_stream_empty;
reg            in_stream_full;
reg     [71:0] slice_stream_buff_0;
reg     [71:0] slice_stream_buff_1;
reg            slice_stream_empty;
reg            slice_stream_full;
reg    [647:0] stencil_stream_buff_0;
reg    [647:0] stencil_stream_buff_1;
reg            stencil_stream_empty;
reg            stencil_stream_full;
wire            arg_0_TREADY;
wire      [7:0] arg_1_TDATA;
wire            arg_1_TVALID;
wire            n0;
wire            n1;
wire            n2;
wire            n3;
wire            n4;
wire            n5;
wire            n6;
wire            n7;
wire            n8;
wire            n9;
wire      [7:0] n10;
wire      [7:0] n11;
wire      [7:0] n12;
wire      [7:0] n13;
wire            n14;
wire            n15;
wire            n16;
wire            n17;
wire            n18;
wire            n19;
wire            n20;
wire            n21;
wire            n22;
wire            n23;
wire            n24;
wire            n25;
wire            n26;
wire            n27;
wire            n28;
wire            n29;
wire            n30;
wire            n31;
wire            n32;
wire            n33;
wire            n34;
wire            n35;
wire            n36;
wire            n37;
wire            n38;
wire            n39;
wire            n40;
wire            n41;
wire            n42;
wire            n43;
wire            n44;
wire     [18:0] n45;
wire     [18:0] n46;
wire            n47;
wire     [18:0] n48;
wire     [18:0] n49;
wire     [18:0] n50;
wire     [18:0] n51;
wire     [18:0] n52;
wire     [18:0] n53;
wire     [18:0] n54;
wire     [18:0] n55;
wire            n56;
wire            n57;
wire     [63:0] n58;
wire     [63:0] n59;
wire     [63:0] n60;
wire     [63:0] n61;
wire     [63:0] n62;
wire     [63:0] n63;
wire     [63:0] n64;
wire     [63:0] n65;
wire     [63:0] n66;
wire            n67;
wire            n68;
wire            n69;
wire      [8:0] n70;
wire      [8:0] n71;
wire      [8:0] n72;
wire      [8:0] n73;
wire      [8:0] n74;
wire      [8:0] n75;
wire      [8:0] n76;
wire      [8:0] n77;
wire            n78;
wire      [9:0] n79;
wire      [9:0] n80;
wire      [9:0] n81;
wire      [9:0] n82;
wire      [9:0] n83;
wire      [9:0] n84;
wire      [9:0] n85;
wire            n86;
wire     [71:0] n87;
wire     [71:0] n88;
wire     [71:0] n89;
wire     [71:0] n90;
wire     [71:0] n91;
wire     [71:0] n92;
wire     [71:0] n93;
wire     [71:0] n94;
wire     [71:0] n95;
wire     [71:0] n96;
wire     [71:0] n97;
wire     [71:0] n98;
wire     [71:0] n99;
wire     [71:0] n100;
wire     [71:0] n101;
wire     [71:0] n102;
wire     [71:0] n103;
wire     [71:0] n104;
wire     [71:0] n105;
wire     [71:0] n106;
wire     [71:0] n107;
wire     [71:0] n108;
wire     [71:0] n109;
wire     [71:0] n110;
wire     [71:0] n111;
wire     [71:0] n112;
wire     [71:0] n113;
wire     [71:0] n114;
wire     [71:0] n115;
wire     [71:0] n116;
wire     [71:0] n117;
wire     [71:0] n118;
wire     [71:0] n119;
wire     [71:0] n120;
wire     [71:0] n121;
wire     [71:0] n122;
wire     [71:0] n123;
wire     [71:0] n124;
wire     [71:0] n125;
wire     [71:0] n126;
wire     [71:0] n127;
wire     [71:0] n128;
wire     [71:0] n129;
wire     [71:0] n130;
wire     [71:0] n131;
wire     [71:0] n132;
wire     [71:0] n133;
wire     [71:0] n134;
wire     [71:0] n135;
wire      [8:0] n136;
wire      [8:0] n137;
wire      [8:0] n138;
wire      [8:0] n139;
wire      [8:0] n140;
wire      [8:0] n141;
wire      [8:0] n142;
wire            n143;
wire            n144;
wire      [9:0] n145;
wire      [9:0] n146;
wire      [9:0] n147;
wire      [9:0] n148;
wire      [9:0] n149;
wire      [9:0] n150;
wire      [9:0] n151;
wire      [9:0] n152;
wire      [9:0] n153;
wire            n154;
wire    [647:0] n155;
wire      [7:0] n156;
wire      [7:0] n157;
wire      [7:0] n158;
wire      [7:0] n159;
wire      [7:0] n160;
wire      [7:0] n161;
wire      [7:0] n162;
wire            n163;
wire            n164;
wire            n165;
wire            n166;
wire            n167;
wire            n168;
wire            n169;
wire            n170;
wire            n171;
wire            n172;
wire            n173;
wire            n174;
wire            n175;
wire            n176;
wire            n177;
wire     [18:0] n178;
wire            n179;
wire            n180;
wire            n181;
wire            n182;
wire            n183;
wire            n184;
wire            n185;
wire            n186;
wire            n187;
wire            n188;
wire            n189;
wire            n190;
wire            n191;
wire            n192;
wire            n193;
wire            n194;
wire            n195;
wire            n196;
wire            n197;
wire            n198;
wire            n199;
wire            n200;
wire            n201;
wire            n202;
wire            n203;
wire            n204;
wire            n205;
wire            n206;
wire            n207;
wire            n208;
wire            n209;
wire            n210;
wire            n211;
wire            n212;
wire            n213;
wire            n214;
wire            n215;
wire            n216;
wire            n217;
wire            n218;
wire            n219;
wire            n220;
wire            n221;
wire            n222;
wire            n223;
wire            n224;
wire            n225;
wire            n226;
wire            n227;
wire            n228;
wire            n229;
wire     [18:0] n230;
wire     [18:0] n231;
wire     [18:0] n232;
wire     [18:0] n233;
wire     [18:0] n234;
wire     [18:0] n235;
wire     [18:0] n236;
wire            n237;
wire            n238;
wire            n239;
wire            n240;
wire            n241;
wire            n242;
wire            n243;
wire            n244;
wire            n245;
wire            n246;
wire            n247;
wire            n248;
wire            n249;
wire            n250;
wire            n251;
wire            n252;
wire            n253;
wire            n254;
wire            n255;
wire            n256;
wire            n257;
wire            n258;
wire            n259;
wire            n260;
wire            n261;
wire            n262;
wire            n263;
wire            n264;
wire            n265;
wire            n266;
wire            n267;
wire            n268;
wire            n269;
wire            n270;
wire            n271;
wire            n272;
wire            n273;
wire            n274;
wire            n275;
wire            n276;
wire            n277;
wire            n278;
wire            n279;
wire            n280;
wire            n281;
wire            n282;
wire            n283;
wire            n284;
wire            n285;
wire            n286;
wire            n287;
wire            n288;
wire            n289;
wire            n290;
wire      [7:0] n291;
wire      [7:0] n292;
wire      [7:0] n293;
wire      [7:0] n294;
wire      [7:0] n295;
wire      [7:0] n296;
wire      [7:0] n297;
wire      [7:0] n298;
wire      [7:0] n299;
wire      [7:0] n300;
wire      [7:0] n301;
wire      [7:0] n302;
wire            n303;
wire            n304;
wire            n305;
wire            n306;
wire            n307;
wire            n308;
wire            n309;
wire            n310;
wire            n311;
wire            n312;
wire            n313;
wire            n314;
wire            n315;
wire            n316;
wire            n317;
wire            n318;
wire      [7:0] n319;
wire            n320;
wire      [7:0] n321;
wire            n322;
wire      [7:0] n323;
wire            n324;
wire      [7:0] n325;
wire            n326;
wire      [7:0] n327;
wire            n328;
wire      [7:0] n329;
wire            n330;
wire      [7:0] n331;
wire            n332;
wire      [7:0] n333;
wire      [7:0] n334;
wire      [7:0] n335;
wire      [7:0] n336;
wire      [7:0] n337;
wire      [7:0] n338;
wire      [7:0] n339;
wire      [7:0] n340;
wire      [7:0] n341;
wire      [7:0] n342;
wire      [7:0] n343;
wire      [7:0] n344;
wire      [7:0] n345;
wire      [7:0] n346;
wire      [7:0] n347;
wire      [7:0] n348;
wire      [7:0] n349;
wire      [7:0] n350;
wire      [7:0] n351;
wire      [7:0] n352;
wire      [7:0] n353;
wire      [7:0] n354;
wire      [7:0] n355;
wire      [7:0] n356;
wire      [7:0] n357;
wire      [7:0] n358;
wire      [7:0] n359;
wire      [7:0] n360;
wire      [7:0] n361;
wire      [7:0] n362;
wire      [7:0] n363;
wire      [7:0] n364;
wire      [7:0] n365;
wire      [7:0] n366;
wire      [7:0] n367;
wire      [7:0] n368;
wire      [7:0] n369;
wire      [7:0] n370;
wire      [7:0] n371;
wire      [7:0] n372;
wire      [7:0] n373;
wire      [7:0] n374;
wire      [7:0] n375;
wire      [7:0] n376;
wire      [7:0] n377;
wire      [7:0] n378;
wire      [7:0] n379;
wire      [7:0] n380;
wire      [7:0] n381;
wire      [7:0] n382;
wire      [7:0] n383;
wire      [7:0] n384;
wire      [7:0] n385;
wire      [7:0] n386;
wire      [7:0] n387;
wire      [7:0] n388;
wire      [7:0] n389;
wire      [7:0] n390;
wire     [15:0] n391;
wire     [23:0] n392;
wire     [31:0] n393;
wire     [39:0] n394;
wire     [47:0] n395;
wire     [55:0] n396;
wire     [63:0] n397;
wire     [71:0] n398;
wire     [71:0] n399;
wire     [71:0] n400;
wire     [71:0] n401;
wire     [71:0] n402;
wire     [71:0] n403;
wire     [71:0] n404;
wire     [71:0] n405;
wire     [71:0] n406;
wire     [71:0] n407;
wire     [71:0] n408;
wire     [71:0] n409;
wire     [71:0] n410;
wire     [71:0] n411;
wire     [71:0] n412;
wire            n413;
wire            n414;
wire            n415;
wire            n416;
wire            n417;
wire            n418;
wire            n419;
wire            n420;
wire            n421;
wire            n422;
wire            n423;
wire            n424;
wire            n425;
wire            n426;
wire            n427;
wire            n428;
wire            n429;
wire            n430;
wire      [7:0] n431;
wire      [7:0] n432;
wire      [7:0] n433;
wire      [7:0] n434;
wire      [7:0] n435;
wire      [7:0] n436;
wire      [7:0] n437;
wire      [7:0] n438;
wire      [7:0] n439;
wire     [15:0] n440;
wire     [23:0] n441;
wire     [31:0] n442;
wire     [39:0] n443;
wire     [47:0] n444;
wire     [55:0] n445;
wire     [63:0] n446;
wire     [71:0] n447;
wire      [7:0] n448;
wire      [7:0] n449;
wire      [7:0] n450;
wire      [7:0] n451;
wire      [7:0] n452;
wire      [7:0] n453;
wire      [7:0] n454;
wire      [7:0] n455;
wire      [7:0] n456;
wire     [15:0] n457;
wire     [23:0] n458;
wire     [31:0] n459;
wire     [39:0] n460;
wire     [47:0] n461;
wire     [55:0] n462;
wire     [63:0] n463;
wire     [71:0] n464;
wire      [7:0] n465;
wire      [7:0] n466;
wire      [7:0] n467;
wire      [7:0] n468;
wire      [7:0] n469;
wire      [7:0] n470;
wire      [7:0] n471;
wire      [7:0] n472;
wire      [7:0] n473;
wire     [15:0] n474;
wire     [23:0] n475;
wire     [31:0] n476;
wire     [39:0] n477;
wire     [47:0] n478;
wire     [55:0] n479;
wire     [63:0] n480;
wire     [71:0] n481;
wire      [7:0] n482;
wire      [7:0] n483;
wire      [7:0] n484;
wire      [7:0] n485;
wire      [7:0] n486;
wire      [7:0] n487;
wire      [7:0] n488;
wire      [7:0] n489;
wire      [7:0] n490;
wire     [15:0] n491;
wire     [23:0] n492;
wire     [31:0] n493;
wire     [39:0] n494;
wire     [47:0] n495;
wire     [55:0] n496;
wire     [63:0] n497;
wire     [71:0] n498;
wire      [7:0] n499;
wire      [7:0] n500;
wire      [7:0] n501;
wire      [7:0] n502;
wire      [7:0] n503;
wire      [7:0] n504;
wire      [7:0] n505;
wire      [7:0] n506;
wire      [7:0] n507;
wire     [15:0] n508;
wire     [23:0] n509;
wire     [31:0] n510;
wire     [39:0] n511;
wire     [47:0] n512;
wire     [55:0] n513;
wire     [63:0] n514;
wire     [71:0] n515;
wire      [7:0] n516;
wire      [7:0] n517;
wire      [7:0] n518;
wire      [7:0] n519;
wire      [7:0] n520;
wire      [7:0] n521;
wire      [7:0] n522;
wire      [7:0] n523;
wire      [7:0] n524;
wire     [15:0] n525;
wire     [23:0] n526;
wire     [31:0] n527;
wire     [39:0] n528;
wire     [47:0] n529;
wire     [55:0] n530;
wire     [63:0] n531;
wire     [71:0] n532;
wire      [7:0] n533;
wire      [7:0] n534;
wire      [7:0] n535;
wire      [7:0] n536;
wire      [7:0] n537;
wire      [7:0] n538;
wire      [7:0] n539;
wire      [7:0] n540;
wire      [7:0] n541;
wire     [15:0] n542;
wire     [23:0] n543;
wire     [31:0] n544;
wire     [39:0] n545;
wire     [47:0] n546;
wire     [55:0] n547;
wire     [63:0] n548;
wire     [71:0] n549;
wire      [7:0] n550;
wire      [7:0] n551;
wire      [7:0] n552;
wire      [7:0] n553;
wire      [7:0] n554;
wire      [7:0] n555;
wire      [7:0] n556;
wire      [7:0] n557;
wire      [7:0] n558;
wire     [15:0] n559;
wire     [23:0] n560;
wire     [31:0] n561;
wire     [39:0] n562;
wire     [47:0] n563;
wire     [55:0] n564;
wire     [63:0] n565;
wire     [71:0] n566;
wire      [7:0] n567;
wire      [7:0] n568;
wire      [7:0] n569;
wire      [7:0] n570;
wire      [7:0] n571;
wire      [7:0] n572;
wire      [7:0] n573;
wire      [7:0] n574;
wire      [7:0] n575;
wire     [15:0] n576;
wire     [23:0] n577;
wire     [31:0] n578;
wire     [39:0] n579;
wire     [47:0] n580;
wire     [55:0] n581;
wire     [63:0] n582;
wire     [71:0] n583;
wire    [143:0] n584;
wire    [215:0] n585;
wire    [287:0] n586;
wire    [359:0] n587;
wire    [431:0] n588;
wire    [503:0] n589;
wire    [575:0] n590;
wire    [647:0] n591;
wire    [647:0] n592;
wire    [647:0] n593;
wire    [647:0] n594;
wire    [647:0] n595;
wire    [647:0] n596;
wire    [647:0] n597;
wire    [647:0] n598;
wire    [647:0] n599;
wire    [647:0] n600;
wire    [647:0] n601;
wire    [647:0] n602;
wire    [647:0] n603;
wire    [647:0] n604;
wire            n605;
wire            n606;
wire            n607;
wire            n608;
wire            n609;
wire            n610;
wire            n611;
wire            n612;
wire            n613;
wire            n614;
wire            n615;
wire            n616;
wire            n617;
wire            n618;
wire            n619;
wire            n620;
wire            n621;
wire            n622;
wire      [8:0] LB2D_proc_0_addr0;
wire      [7:0] LB2D_proc_0_data0;
wire            n623;
wire            n624;
wire            n625;
wire            n626;
wire            n627;
wire            n628;
wire            n629;
wire            n630;
wire            n631;
wire            n632;
wire            n633;
wire            n634;
wire            n635;
wire            n636;
wire            n637;
wire            n638;
wire            n639;
wire            n640;
wire            n641;
wire      [8:0] LB2D_proc_1_addr0;
wire      [7:0] LB2D_proc_1_data0;
wire            n642;
wire            n643;
wire            n644;
wire      [8:0] LB2D_proc_2_addr0;
wire      [7:0] LB2D_proc_2_data0;
wire            n645;
wire            n646;
wire            n647;
wire      [8:0] LB2D_proc_3_addr0;
wire      [7:0] LB2D_proc_3_data0;
wire            n648;
wire            n649;
wire            n650;
wire      [8:0] LB2D_proc_4_addr0;
wire      [7:0] LB2D_proc_4_data0;
wire            n651;
wire            n652;
wire            n653;
wire      [8:0] LB2D_proc_5_addr0;
wire      [7:0] LB2D_proc_5_data0;
wire            n654;
wire            n655;
wire            n656;
wire      [8:0] LB2D_proc_6_addr0;
wire      [7:0] LB2D_proc_6_data0;
wire            n657;
wire            n658;
wire            n659;
wire      [8:0] LB2D_proc_7_addr0;
wire      [7:0] LB2D_proc_7_data0;
wire            n660;
wire            n661;
wire            n662;
wire            n663;
reg      [7:0] LB2D_proc_0[511:0];
reg      [7:0] LB2D_proc_1[511:0];
reg      [7:0] LB2D_proc_2[511:0];
reg      [7:0] LB2D_proc_3[511:0];
reg      [7:0] LB2D_proc_4[511:0];
reg      [7:0] LB2D_proc_5[511:0];
reg      [7:0] LB2D_proc_6[511:0];
reg      [7:0] LB2D_proc_7[511:0];
wire clk;
wire rst;
wire step;
assign n0 =  ( arg_1_TREADY ) == ( 1'd1 )  ;
assign n1 =  ( arg_1_TVALID ) == ( 1'd1 )  ;
assign n2 =  ( n0 ) & ( n1 )  ;
assign n3 =  ( arg_0_TREADY ) == ( 1'd0 )  ;
assign n4 =  ( n2 ) & ( n3 )  ;
assign n5 =  ( arg_1_TREADY ) == ( 1'd0 )  ;
assign n6 =  ( in_stream_full ) == ( 1'd0 )  ;
assign n7 =  ( n5 ) & ( n6 )  ;
assign n8 =  ( LB1D_it_1 ) == ( 1'd1 )  ;
assign n9 =  ( n7 ) & ( n8 )  ;
assign n10 =  ( n9 ) ? ( LB1D_in ) : ( LB1D_buff ) ;
assign n11 =  ( n4 ) ? ( LB1D_buff ) : ( n10 ) ;
assign n12 =  ( n9 ) ? ( arg_1_TDATA ) : ( LB1D_in ) ;
assign n13 =  ( n4 ) ? ( LB1D_in ) : ( n12 ) ;
assign n14 =  ( LB1D_it_1 ) == ( 1'd0 )  ;
assign n15 =  ( n7 ) & ( n14 )  ;
assign n16 =  ( n15 ) ? ( 1'd1 ) : ( LB1D_it_1 ) ;
assign n17 =  ( arg_0_TREADY ) == ( 1'd1 )  ;
assign n18 =  ( arg_0_TVALID ) == ( 1'd1 )  ;
assign n19 =  ( n17 ) & ( n18 )  ;
assign n20 =  ( arg_1_TVALID ) == ( 1'd0 )  ;
assign n21 =  ( n19 ) & ( n20 )  ;
assign n22 =  ( arg_0_TVALID ) == ( 1'd0 )  ;
assign n23 =  ( gb_exit_it_1 ) == ( 1'd0 )  ;
assign n24 =  ( stencil_stream_empty ) == ( 1'd0 )  ;
assign n25 =  ( n23 ) & ( n24 )  ;
assign n26 =  ( gb_exit_it_1 ) == ( 1'd1 )  ;
assign n27 =  ( gb_exit_it_8 ) == ( 1'd0 )  ;
assign n28 =  ( n26 ) & ( n27 )  ;
assign n29 =  ( n25 ) | ( n28 )  ;
assign n30 =  ( n22 ) & ( n29 )  ;
assign n31 =  ( slice_stream_empty ) == ( 1'd0 )  ;
assign n32 =  ( LB2D_shift_x ) != ( 9'd488 )  ;
assign n33 =  ( n31 ) & ( n32 )  ;
assign n34 =  ( stencil_stream_full ) == ( 1'd0 )  ;
assign n35 =  ( LB2D_shift_x ) < ( 9'd8 )  ;
assign n36 =  ( n34 ) | ( n35 )  ;
assign n37 =  ( n33 ) & ( n36 )  ;
assign n38 =  ( in_stream_empty ) == ( 1'd0 )  ;
assign n39 =  ( LB2D_proc_x ) != ( 9'd488 )  ;
assign n40 =  ( n38 ) & ( n39 )  ;
assign n41 =  ( slice_stream_full ) == ( 1'd0 )  ;
assign n42 =  ( LB2D_proc_y ) < ( 10'd8 )  ;
assign n43 =  ( n41 ) | ( n42 )  ;
assign n44 =  ( n40 ) & ( n43 )  ;
assign n45 =  ( LB1D_p_cnt ) + ( 19'd1 )  ;
assign n46 =  ( 19'd316224 ) - ( 19'd1 )  ;
assign n47 =  ( LB1D_p_cnt ) == ( n46 )  ;
assign n48 =  ( n47 ) ? ( 19'd0 ) : ( n45 ) ;
assign n49 =  ( n9 ) ? ( n48 ) : ( LB1D_p_cnt ) ;
assign n50 =  ( n15 ) ? ( n45 ) : ( n49 ) ;
assign n51 =  ( n44 ) ? ( LB1D_p_cnt ) : ( n50 ) ;
assign n52 =  ( n37 ) ? ( LB1D_p_cnt ) : ( n51 ) ;
assign n53 =  ( n30 ) ? ( LB1D_p_cnt ) : ( n52 ) ;
assign n54 =  ( n4 ) ? ( LB1D_p_cnt ) : ( n53 ) ;
assign n55 =  ( n21 ) ? ( LB1D_p_cnt ) : ( n54 ) ;
assign n56 =  ( LB2D_proc_w ) < ( 64'd7 )  ;
assign n57 =  ( LB2D_proc_x ) < ( 9'd488 )  ;
assign n58 =  ( LB2D_proc_w ) + ( 64'd1 )  ;
assign n59 =  ( n57 ) ? ( LB2D_proc_w ) : ( n58 ) ;
assign n60 =  ( n56 ) ? ( n59 ) : ( 64'd0 ) ;
assign n61 =  ( n9 ) ? ( LB2D_proc_w ) : ( LB2D_proc_w ) ;
assign n62 =  ( n44 ) ? ( n60 ) : ( n61 ) ;
assign n63 =  ( n37 ) ? ( LB2D_proc_w ) : ( n62 ) ;
assign n64 =  ( n30 ) ? ( LB2D_proc_w ) : ( n63 ) ;
assign n65 =  ( n4 ) ? ( LB2D_proc_w ) : ( n64 ) ;
assign n66 =  ( n21 ) ? ( LB2D_proc_w ) : ( n65 ) ;
assign n67 =  ( LB2D_proc_x ) == ( 9'd488 )  ;
assign n68 =  ( n38 ) & ( n67 )  ;
assign n69 =  ( n68 ) & ( n43 )  ;
assign n70 =  ( LB2D_proc_x ) + ( 9'd1 )  ;
assign n71 =  ( n9 ) ? ( LB2D_proc_x ) : ( LB2D_proc_x ) ;
assign n72 =  ( n44 ) ? ( n70 ) : ( n71 ) ;
assign n73 =  ( n69 ) ? ( 9'd0 ) : ( n72 ) ;
assign n74 =  ( n37 ) ? ( LB2D_proc_x ) : ( n73 ) ;
assign n75 =  ( n30 ) ? ( LB2D_proc_x ) : ( n74 ) ;
assign n76 =  ( n4 ) ? ( LB2D_proc_x ) : ( n75 ) ;
assign n77 =  ( n21 ) ? ( LB2D_proc_x ) : ( n76 ) ;
assign n78 =  ( LB2D_proc_y ) < ( 10'd488 )  ;
assign n79 =  ( n78 ) ? ( LB2D_proc_y ) : ( 10'd488 ) ;
assign n80 =  ( n9 ) ? ( LB2D_proc_y ) : ( LB2D_proc_y ) ;
assign n81 =  ( n44 ) ? ( n79 ) : ( n80 ) ;
assign n82 =  ( n37 ) ? ( LB2D_proc_y ) : ( n81 ) ;
assign n83 =  ( n30 ) ? ( LB2D_proc_y ) : ( n82 ) ;
assign n84 =  ( n4 ) ? ( LB2D_proc_y ) : ( n83 ) ;
assign n85 =  ( n21 ) ? ( LB2D_proc_y ) : ( n84 ) ;
assign n86 =  ( slice_stream_full ) == ( 1'd1 )  ;
assign n87 =  ( n86 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n88 =  ( n9 ) ? ( LB2D_shift_0 ) : ( LB2D_shift_0 ) ;
assign n89 =  ( n44 ) ? ( LB2D_shift_0 ) : ( n88 ) ;
assign n90 =  ( n37 ) ? ( n87 ) : ( n89 ) ;
assign n91 =  ( n30 ) ? ( LB2D_shift_0 ) : ( n90 ) ;
assign n92 =  ( n4 ) ? ( LB2D_shift_0 ) : ( n91 ) ;
assign n93 =  ( n21 ) ? ( LB2D_shift_0 ) : ( n92 ) ;
assign n94 =  ( n9 ) ? ( LB2D_shift_1 ) : ( LB2D_shift_1 ) ;
assign n95 =  ( n44 ) ? ( LB2D_shift_1 ) : ( n94 ) ;
assign n96 =  ( n37 ) ? ( LB2D_shift_0 ) : ( n95 ) ;
assign n97 =  ( n30 ) ? ( LB2D_shift_1 ) : ( n96 ) ;
assign n98 =  ( n4 ) ? ( LB2D_shift_1 ) : ( n97 ) ;
assign n99 =  ( n21 ) ? ( LB2D_shift_1 ) : ( n98 ) ;
assign n100 =  ( n9 ) ? ( LB2D_shift_2 ) : ( LB2D_shift_2 ) ;
assign n101 =  ( n44 ) ? ( LB2D_shift_2 ) : ( n100 ) ;
assign n102 =  ( n37 ) ? ( LB2D_shift_1 ) : ( n101 ) ;
assign n103 =  ( n30 ) ? ( LB2D_shift_2 ) : ( n102 ) ;
assign n104 =  ( n4 ) ? ( LB2D_shift_2 ) : ( n103 ) ;
assign n105 =  ( n21 ) ? ( LB2D_shift_2 ) : ( n104 ) ;
assign n106 =  ( n9 ) ? ( LB2D_shift_3 ) : ( LB2D_shift_3 ) ;
assign n107 =  ( n44 ) ? ( LB2D_shift_3 ) : ( n106 ) ;
assign n108 =  ( n37 ) ? ( LB2D_shift_2 ) : ( n107 ) ;
assign n109 =  ( n30 ) ? ( LB2D_shift_3 ) : ( n108 ) ;
assign n110 =  ( n4 ) ? ( LB2D_shift_3 ) : ( n109 ) ;
assign n111 =  ( n21 ) ? ( LB2D_shift_3 ) : ( n110 ) ;
assign n112 =  ( n9 ) ? ( LB2D_shift_4 ) : ( LB2D_shift_4 ) ;
assign n113 =  ( n44 ) ? ( LB2D_shift_4 ) : ( n112 ) ;
assign n114 =  ( n37 ) ? ( LB2D_shift_3 ) : ( n113 ) ;
assign n115 =  ( n30 ) ? ( LB2D_shift_4 ) : ( n114 ) ;
assign n116 =  ( n4 ) ? ( LB2D_shift_4 ) : ( n115 ) ;
assign n117 =  ( n21 ) ? ( LB2D_shift_4 ) : ( n116 ) ;
assign n118 =  ( n9 ) ? ( LB2D_shift_5 ) : ( LB2D_shift_5 ) ;
assign n119 =  ( n44 ) ? ( LB2D_shift_5 ) : ( n118 ) ;
assign n120 =  ( n37 ) ? ( LB2D_shift_4 ) : ( n119 ) ;
assign n121 =  ( n30 ) ? ( LB2D_shift_5 ) : ( n120 ) ;
assign n122 =  ( n4 ) ? ( LB2D_shift_5 ) : ( n121 ) ;
assign n123 =  ( n21 ) ? ( LB2D_shift_5 ) : ( n122 ) ;
assign n124 =  ( n9 ) ? ( LB2D_shift_6 ) : ( LB2D_shift_6 ) ;
assign n125 =  ( n44 ) ? ( LB2D_shift_6 ) : ( n124 ) ;
assign n126 =  ( n37 ) ? ( LB2D_shift_5 ) : ( n125 ) ;
assign n127 =  ( n30 ) ? ( LB2D_shift_6 ) : ( n126 ) ;
assign n128 =  ( n4 ) ? ( LB2D_shift_6 ) : ( n127 ) ;
assign n129 =  ( n21 ) ? ( LB2D_shift_6 ) : ( n128 ) ;
assign n130 =  ( n9 ) ? ( LB2D_shift_7 ) : ( LB2D_shift_7 ) ;
assign n131 =  ( n44 ) ? ( LB2D_shift_7 ) : ( n130 ) ;
assign n132 =  ( n37 ) ? ( LB2D_shift_6 ) : ( n131 ) ;
assign n133 =  ( n30 ) ? ( LB2D_shift_7 ) : ( n132 ) ;
assign n134 =  ( n4 ) ? ( LB2D_shift_7 ) : ( n133 ) ;
assign n135 =  ( n21 ) ? ( LB2D_shift_7 ) : ( n134 ) ;
assign n136 =  ( LB2D_shift_x ) + ( 9'd1 )  ;
assign n137 =  ( n9 ) ? ( LB2D_shift_x ) : ( LB2D_shift_x ) ;
assign n138 =  ( n44 ) ? ( LB2D_shift_x ) : ( n137 ) ;
assign n139 =  ( n37 ) ? ( n136 ) : ( n138 ) ;
assign n140 =  ( n30 ) ? ( LB2D_shift_x ) : ( n139 ) ;
assign n141 =  ( n4 ) ? ( LB2D_shift_x ) : ( n140 ) ;
assign n142 =  ( n21 ) ? ( LB2D_shift_x ) : ( n141 ) ;
assign n143 =  ( LB2D_shift_y ) < ( 10'd480 )  ;
assign n144 =  ( LB2D_shift_x ) < ( 9'd488 )  ;
assign n145 =  ( LB2D_shift_y ) + ( 10'd1 )  ;
assign n146 =  ( n144 ) ? ( LB2D_shift_y ) : ( n145 ) ;
assign n147 =  ( n143 ) ? ( n146 ) : ( 10'd480 ) ;
assign n148 =  ( n9 ) ? ( LB2D_shift_y ) : ( LB2D_shift_y ) ;
assign n149 =  ( n44 ) ? ( LB2D_shift_y ) : ( n148 ) ;
assign n150 =  ( n37 ) ? ( n147 ) : ( n149 ) ;
assign n151 =  ( n30 ) ? ( LB2D_shift_y ) : ( n150 ) ;
assign n152 =  ( n4 ) ? ( LB2D_shift_y ) : ( n151 ) ;
assign n153 =  ( n21 ) ? ( LB2D_shift_y ) : ( n152 ) ;
assign n154 =  ( stencil_stream_full ) == ( 1'd1 )  ;
assign n155 =  ( n154 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_0 ) ;
//assign n156 = gb_fun(n155) ;
gb_fun gb_fun_U (
        .stencil (n155),
        .res (n156)
        );
assign n157 =  ( n9 ) ? ( arg_0_TDATA ) : ( arg_0_TDATA ) ;
assign n158 =  ( n44 ) ? ( arg_0_TDATA ) : ( n157 ) ;
assign n159 =  ( n37 ) ? ( arg_0_TDATA ) : ( n158 ) ;
assign n160 =  ( n30 ) ? ( n156 ) : ( n159 ) ;
assign n161 =  ( n4 ) ? ( arg_0_TDATA ) : ( n160 ) ;
assign n162 =  ( n21 ) ? ( arg_0_TDATA ) : ( n161 ) ;
assign n163 =  ( gb_pp_it_8 ) == ( 1'd1 )  ;
assign n164 =  ( n163 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n165 =  ( n9 ) ? ( arg_0_TVALID ) : ( arg_0_TVALID ) ;
assign n166 =  ( n44 ) ? ( arg_0_TVALID ) : ( n165 ) ;
assign n167 =  ( n37 ) ? ( arg_0_TVALID ) : ( n166 ) ;
assign n168 =  ( n30 ) ? ( n164 ) : ( n167 ) ;
assign n169 =  ( n4 ) ? ( arg_0_TVALID ) : ( n168 ) ;
assign n170 =  ( n21 ) ? ( 1'd0 ) : ( n169 ) ;
assign n171 =  ( n9 ) ? ( 1'd1 ) : ( arg_1_TREADY ) ;
assign n172 =  ( n15 ) ? ( 1'd1 ) : ( n171 ) ;
assign n173 =  ( n44 ) ? ( arg_1_TREADY ) : ( n172 ) ;
assign n174 =  ( n37 ) ? ( arg_1_TREADY ) : ( n173 ) ;
assign n175 =  ( n30 ) ? ( arg_1_TREADY ) : ( n174 ) ;
assign n176 =  ( n4 ) ? ( 1'd0 ) : ( n175 ) ;
assign n177 =  ( n21 ) ? ( 1'd0 ) : ( n176 ) ;
assign n178 =  ( gb_p_cnt ) + ( 19'd1 )  ;
assign n179 =  ( n178 ) == ( 19'd307200 )  ;
assign n180 =  ( n179 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n181 =  ( n9 ) ? ( gb_exit_it_1 ) : ( gb_exit_it_1 ) ;
assign n182 =  ( n44 ) ? ( gb_exit_it_1 ) : ( n181 ) ;
assign n183 =  ( n37 ) ? ( gb_exit_it_1 ) : ( n182 ) ;
assign n184 =  ( n30 ) ? ( n180 ) : ( n183 ) ;
assign n185 =  ( n4 ) ? ( gb_exit_it_1 ) : ( n184 ) ;
assign n186 =  ( n21 ) ? ( gb_exit_it_1 ) : ( n185 ) ;
assign n187 =  ( n9 ) ? ( gb_exit_it_2 ) : ( gb_exit_it_2 ) ;
assign n188 =  ( n44 ) ? ( gb_exit_it_2 ) : ( n187 ) ;
assign n189 =  ( n37 ) ? ( gb_exit_it_2 ) : ( n188 ) ;
assign n190 =  ( n30 ) ? ( gb_exit_it_1 ) : ( n189 ) ;
assign n191 =  ( n4 ) ? ( gb_exit_it_2 ) : ( n190 ) ;
assign n192 =  ( n21 ) ? ( gb_exit_it_2 ) : ( n191 ) ;
assign n193 =  ( n9 ) ? ( gb_exit_it_3 ) : ( gb_exit_it_3 ) ;
assign n194 =  ( n44 ) ? ( gb_exit_it_3 ) : ( n193 ) ;
assign n195 =  ( n37 ) ? ( gb_exit_it_3 ) : ( n194 ) ;
assign n196 =  ( n30 ) ? ( gb_exit_it_2 ) : ( n195 ) ;
assign n197 =  ( n4 ) ? ( gb_exit_it_3 ) : ( n196 ) ;
assign n198 =  ( n21 ) ? ( gb_exit_it_3 ) : ( n197 ) ;
assign n199 =  ( n9 ) ? ( gb_exit_it_4 ) : ( gb_exit_it_4 ) ;
assign n200 =  ( n44 ) ? ( gb_exit_it_4 ) : ( n199 ) ;
assign n201 =  ( n37 ) ? ( gb_exit_it_4 ) : ( n200 ) ;
assign n202 =  ( n30 ) ? ( gb_exit_it_3 ) : ( n201 ) ;
assign n203 =  ( n4 ) ? ( gb_exit_it_4 ) : ( n202 ) ;
assign n204 =  ( n21 ) ? ( gb_exit_it_4 ) : ( n203 ) ;
assign n205 =  ( n9 ) ? ( gb_exit_it_5 ) : ( gb_exit_it_5 ) ;
assign n206 =  ( n44 ) ? ( gb_exit_it_5 ) : ( n205 ) ;
assign n207 =  ( n37 ) ? ( gb_exit_it_5 ) : ( n206 ) ;
assign n208 =  ( n30 ) ? ( gb_exit_it_4 ) : ( n207 ) ;
assign n209 =  ( n4 ) ? ( gb_exit_it_5 ) : ( n208 ) ;
assign n210 =  ( n21 ) ? ( gb_exit_it_5 ) : ( n209 ) ;
assign n211 =  ( n9 ) ? ( gb_exit_it_6 ) : ( gb_exit_it_6 ) ;
assign n212 =  ( n44 ) ? ( gb_exit_it_6 ) : ( n211 ) ;
assign n213 =  ( n37 ) ? ( gb_exit_it_6 ) : ( n212 ) ;
assign n214 =  ( n30 ) ? ( gb_exit_it_5 ) : ( n213 ) ;
assign n215 =  ( n4 ) ? ( gb_exit_it_6 ) : ( n214 ) ;
assign n216 =  ( n21 ) ? ( gb_exit_it_6 ) : ( n215 ) ;
assign n217 =  ( n9 ) ? ( gb_exit_it_7 ) : ( gb_exit_it_7 ) ;
assign n218 =  ( n44 ) ? ( gb_exit_it_7 ) : ( n217 ) ;
assign n219 =  ( n37 ) ? ( gb_exit_it_7 ) : ( n218 ) ;
assign n220 =  ( n30 ) ? ( gb_exit_it_6 ) : ( n219 ) ;
assign n221 =  ( n4 ) ? ( gb_exit_it_7 ) : ( n220 ) ;
assign n222 =  ( n21 ) ? ( gb_exit_it_7 ) : ( n221 ) ;
assign n223 =  ( n9 ) ? ( gb_exit_it_8 ) : ( gb_exit_it_8 ) ;
assign n224 =  ( n44 ) ? ( gb_exit_it_8 ) : ( n223 ) ;
assign n225 =  ( n37 ) ? ( gb_exit_it_8 ) : ( n224 ) ;
assign n226 =  ( n30 ) ? ( gb_exit_it_7 ) : ( n225 ) ;
assign n227 =  ( n4 ) ? ( gb_exit_it_8 ) : ( n226 ) ;
assign n228 =  ( n21 ) ? ( gb_exit_it_8 ) : ( n227 ) ;
assign n229 =  ( gb_p_cnt ) < ( 19'd307200 )  ;
assign n230 =  ( n229 ) ? ( n178 ) : ( 19'd307200 ) ;
assign n231 =  ( n9 ) ? ( gb_p_cnt ) : ( gb_p_cnt ) ;
assign n232 =  ( n44 ) ? ( gb_p_cnt ) : ( n231 ) ;
assign n233 =  ( n37 ) ? ( gb_p_cnt ) : ( n232 ) ;
assign n234 =  ( n30 ) ? ( n230 ) : ( n233 ) ;
assign n235 =  ( n4 ) ? ( gb_p_cnt ) : ( n234 ) ;
assign n236 =  ( n21 ) ? ( gb_p_cnt ) : ( n235 ) ;
assign n237 =  ( n9 ) ? ( gb_pp_it_1 ) : ( gb_pp_it_1 ) ;
assign n238 =  ( n44 ) ? ( gb_pp_it_1 ) : ( n237 ) ;
assign n239 =  ( n37 ) ? ( gb_pp_it_1 ) : ( n238 ) ;
assign n240 =  ( n30 ) ? ( 1'd1 ) : ( n239 ) ;
assign n241 =  ( n4 ) ? ( gb_pp_it_1 ) : ( n240 ) ;
assign n242 =  ( n21 ) ? ( gb_pp_it_1 ) : ( n241 ) ;
assign n243 =  ( n9 ) ? ( gb_pp_it_2 ) : ( gb_pp_it_2 ) ;
assign n244 =  ( n44 ) ? ( gb_pp_it_2 ) : ( n243 ) ;
assign n245 =  ( n37 ) ? ( gb_pp_it_2 ) : ( n244 ) ;
assign n246 =  ( n30 ) ? ( gb_pp_it_1 ) : ( n245 ) ;
assign n247 =  ( n4 ) ? ( gb_pp_it_2 ) : ( n246 ) ;
assign n248 =  ( n21 ) ? ( gb_pp_it_2 ) : ( n247 ) ;
assign n249 =  ( n9 ) ? ( gb_pp_it_3 ) : ( gb_pp_it_3 ) ;
assign n250 =  ( n44 ) ? ( gb_pp_it_3 ) : ( n249 ) ;
assign n251 =  ( n37 ) ? ( gb_pp_it_3 ) : ( n250 ) ;
assign n252 =  ( n30 ) ? ( gb_pp_it_2 ) : ( n251 ) ;
assign n253 =  ( n4 ) ? ( gb_pp_it_3 ) : ( n252 ) ;
assign n254 =  ( n21 ) ? ( gb_pp_it_3 ) : ( n253 ) ;
assign n255 =  ( n9 ) ? ( gb_pp_it_4 ) : ( gb_pp_it_4 ) ;
assign n256 =  ( n44 ) ? ( gb_pp_it_4 ) : ( n255 ) ;
assign n257 =  ( n37 ) ? ( gb_pp_it_4 ) : ( n256 ) ;
assign n258 =  ( n30 ) ? ( gb_pp_it_3 ) : ( n257 ) ;
assign n259 =  ( n4 ) ? ( gb_pp_it_4 ) : ( n258 ) ;
assign n260 =  ( n21 ) ? ( gb_pp_it_4 ) : ( n259 ) ;
assign n261 =  ( n9 ) ? ( gb_pp_it_5 ) : ( gb_pp_it_5 ) ;
assign n262 =  ( n44 ) ? ( gb_pp_it_5 ) : ( n261 ) ;
assign n263 =  ( n37 ) ? ( gb_pp_it_5 ) : ( n262 ) ;
assign n264 =  ( n30 ) ? ( gb_pp_it_4 ) : ( n263 ) ;
assign n265 =  ( n4 ) ? ( gb_pp_it_5 ) : ( n264 ) ;
assign n266 =  ( n21 ) ? ( gb_pp_it_5 ) : ( n265 ) ;
assign n267 =  ( n9 ) ? ( gb_pp_it_6 ) : ( gb_pp_it_6 ) ;
assign n268 =  ( n44 ) ? ( gb_pp_it_6 ) : ( n267 ) ;
assign n269 =  ( n37 ) ? ( gb_pp_it_6 ) : ( n268 ) ;
assign n270 =  ( n30 ) ? ( gb_pp_it_5 ) : ( n269 ) ;
assign n271 =  ( n4 ) ? ( gb_pp_it_6 ) : ( n270 ) ;
assign n272 =  ( n21 ) ? ( gb_pp_it_6 ) : ( n271 ) ;
assign n273 =  ( n9 ) ? ( gb_pp_it_7 ) : ( gb_pp_it_7 ) ;
assign n274 =  ( n44 ) ? ( gb_pp_it_7 ) : ( n273 ) ;
assign n275 =  ( n37 ) ? ( gb_pp_it_7 ) : ( n274 ) ;
assign n276 =  ( n30 ) ? ( gb_pp_it_6 ) : ( n275 ) ;
assign n277 =  ( n4 ) ? ( gb_pp_it_7 ) : ( n276 ) ;
assign n278 =  ( n21 ) ? ( gb_pp_it_7 ) : ( n277 ) ;
assign n279 =  ( n9 ) ? ( gb_pp_it_8 ) : ( gb_pp_it_8 ) ;
assign n280 =  ( n44 ) ? ( gb_pp_it_8 ) : ( n279 ) ;
assign n281 =  ( n37 ) ? ( gb_pp_it_8 ) : ( n280 ) ;
assign n282 =  ( n30 ) ? ( gb_pp_it_7 ) : ( n281 ) ;
assign n283 =  ( n4 ) ? ( gb_pp_it_8 ) : ( n282 ) ;
assign n284 =  ( n21 ) ? ( gb_pp_it_8 ) : ( n283 ) ;
assign n285 =  ( n9 ) ? ( gb_pp_it_9 ) : ( gb_pp_it_9 ) ;
assign n286 =  ( n44 ) ? ( gb_pp_it_9 ) : ( n285 ) ;
assign n287 =  ( n37 ) ? ( gb_pp_it_9 ) : ( n286 ) ;
assign n288 =  ( n30 ) ? ( gb_pp_it_8 ) : ( n287 ) ;
assign n289 =  ( n4 ) ? ( gb_pp_it_9 ) : ( n288 ) ;
assign n290 =  ( n21 ) ? ( gb_pp_it_9 ) : ( n289 ) ;
assign n291 =  ( n9 ) ? ( LB1D_buff ) : ( in_stream_buff_0 ) ;
assign n292 =  ( n44 ) ? ( in_stream_buff_0 ) : ( n291 ) ;
assign n293 =  ( n37 ) ? ( in_stream_buff_0 ) : ( n292 ) ;
assign n294 =  ( n30 ) ? ( in_stream_buff_0 ) : ( n293 ) ;
assign n295 =  ( n4 ) ? ( in_stream_buff_0 ) : ( n294 ) ;
assign n296 =  ( n21 ) ? ( in_stream_buff_0 ) : ( n295 ) ;
assign n297 =  ( n9 ) ? ( in_stream_buff_0 ) : ( in_stream_buff_1 ) ;
assign n298 =  ( n44 ) ? ( in_stream_buff_1 ) : ( n297 ) ;
assign n299 =  ( n37 ) ? ( in_stream_buff_1 ) : ( n298 ) ;
assign n300 =  ( n30 ) ? ( in_stream_buff_1 ) : ( n299 ) ;
assign n301 =  ( n4 ) ? ( in_stream_buff_1 ) : ( n300 ) ;
assign n302 =  ( n21 ) ? ( in_stream_buff_1 ) : ( n301 ) ;
assign n303 =  ( in_stream_full ) == ( 1'd1 )  ;
assign n304 =  ( n303 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n305 =  ( n9 ) ? ( 1'd0 ) : ( in_stream_empty ) ;
assign n306 =  ( n44 ) ? ( n304 ) : ( n305 ) ;
assign n307 =  ( n37 ) ? ( in_stream_empty ) : ( n306 ) ;
assign n308 =  ( n30 ) ? ( in_stream_empty ) : ( n307 ) ;
assign n309 =  ( n4 ) ? ( in_stream_empty ) : ( n308 ) ;
assign n310 =  ( n21 ) ? ( in_stream_empty ) : ( n309 ) ;
assign n311 =  ( in_stream_empty ) == ( 1'd1 )  ;
assign n312 =  ( n311 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n313 =  ( n9 ) ? ( n312 ) : ( in_stream_full ) ;
assign n314 =  ( n44 ) ? ( 1'd0 ) : ( n313 ) ;
assign n315 =  ( n37 ) ? ( in_stream_full ) : ( n314 ) ;
assign n316 =  ( n30 ) ? ( in_stream_full ) : ( n315 ) ;
assign n317 =  ( n4 ) ? ( in_stream_full ) : ( n316 ) ;
assign n318 =  ( n21 ) ? ( in_stream_full ) : ( n317 ) ;
assign n319 =  ( n303 ) ? ( in_stream_buff_1 ) : ( in_stream_buff_0 ) ;
assign n320 =  ( LB2D_proc_w ) == ( 64'd0 )  ;
assign n321 =  (  LB2D_proc_7 [ LB2D_proc_x ] )  ;
assign n322 =  ( LB2D_proc_w ) == ( 64'd1 )  ;
assign n323 =  (  LB2D_proc_0 [ LB2D_proc_x ] )  ;
assign n324 =  ( LB2D_proc_w ) == ( 64'd2 )  ;
assign n325 =  (  LB2D_proc_1 [ LB2D_proc_x ] )  ;
assign n326 =  ( LB2D_proc_w ) == ( 64'd3 )  ;
assign n327 =  (  LB2D_proc_2 [ LB2D_proc_x ] )  ;
assign n328 =  ( LB2D_proc_w ) == ( 64'd4 )  ;
assign n329 =  (  LB2D_proc_3 [ LB2D_proc_x ] )  ;
assign n330 =  ( LB2D_proc_w ) == ( 64'd5 )  ;
assign n331 =  (  LB2D_proc_4 [ LB2D_proc_x ] )  ;
assign n332 =  ( LB2D_proc_w ) == ( 64'd6 )  ;
assign n333 =  (  LB2D_proc_5 [ LB2D_proc_x ] )  ;
assign n334 =  (  LB2D_proc_6 [ LB2D_proc_x ] )  ;
assign n335 =  ( n332 ) ? ( n333 ) : ( n334 ) ;
assign n336 =  ( n330 ) ? ( n331 ) : ( n335 ) ;
assign n337 =  ( n328 ) ? ( n329 ) : ( n336 ) ;
assign n338 =  ( n326 ) ? ( n327 ) : ( n337 ) ;
assign n339 =  ( n324 ) ? ( n325 ) : ( n338 ) ;
assign n340 =  ( n322 ) ? ( n323 ) : ( n339 ) ;
assign n341 =  ( n320 ) ? ( n321 ) : ( n340 ) ;
assign n342 =  ( n332 ) ? ( n331 ) : ( n333 ) ;
assign n343 =  ( n330 ) ? ( n329 ) : ( n342 ) ;
assign n344 =  ( n328 ) ? ( n327 ) : ( n343 ) ;
assign n345 =  ( n326 ) ? ( n325 ) : ( n344 ) ;
assign n346 =  ( n324 ) ? ( n323 ) : ( n345 ) ;
assign n347 =  ( n322 ) ? ( n321 ) : ( n346 ) ;
assign n348 =  ( n320 ) ? ( n334 ) : ( n347 ) ;
assign n349 =  ( n332 ) ? ( n329 ) : ( n331 ) ;
assign n350 =  ( n330 ) ? ( n327 ) : ( n349 ) ;
assign n351 =  ( n328 ) ? ( n325 ) : ( n350 ) ;
assign n352 =  ( n326 ) ? ( n323 ) : ( n351 ) ;
assign n353 =  ( n324 ) ? ( n321 ) : ( n352 ) ;
assign n354 =  ( n322 ) ? ( n334 ) : ( n353 ) ;
assign n355 =  ( n320 ) ? ( n333 ) : ( n354 ) ;
assign n356 =  ( n332 ) ? ( n327 ) : ( n329 ) ;
assign n357 =  ( n330 ) ? ( n325 ) : ( n356 ) ;
assign n358 =  ( n328 ) ? ( n323 ) : ( n357 ) ;
assign n359 =  ( n326 ) ? ( n321 ) : ( n358 ) ;
assign n360 =  ( n324 ) ? ( n334 ) : ( n359 ) ;
assign n361 =  ( n322 ) ? ( n333 ) : ( n360 ) ;
assign n362 =  ( n320 ) ? ( n331 ) : ( n361 ) ;
assign n363 =  ( n332 ) ? ( n325 ) : ( n327 ) ;
assign n364 =  ( n330 ) ? ( n323 ) : ( n363 ) ;
assign n365 =  ( n328 ) ? ( n321 ) : ( n364 ) ;
assign n366 =  ( n326 ) ? ( n334 ) : ( n365 ) ;
assign n367 =  ( n324 ) ? ( n333 ) : ( n366 ) ;
assign n368 =  ( n322 ) ? ( n331 ) : ( n367 ) ;
assign n369 =  ( n320 ) ? ( n329 ) : ( n368 ) ;
assign n370 =  ( n332 ) ? ( n323 ) : ( n325 ) ;
assign n371 =  ( n330 ) ? ( n321 ) : ( n370 ) ;
assign n372 =  ( n328 ) ? ( n334 ) : ( n371 ) ;
assign n373 =  ( n326 ) ? ( n333 ) : ( n372 ) ;
assign n374 =  ( n324 ) ? ( n331 ) : ( n373 ) ;
assign n375 =  ( n322 ) ? ( n329 ) : ( n374 ) ;
assign n376 =  ( n320 ) ? ( n327 ) : ( n375 ) ;
assign n377 =  ( n332 ) ? ( n321 ) : ( n323 ) ;
assign n378 =  ( n330 ) ? ( n334 ) : ( n377 ) ;
assign n379 =  ( n328 ) ? ( n333 ) : ( n378 ) ;
assign n380 =  ( n326 ) ? ( n331 ) : ( n379 ) ;
assign n381 =  ( n324 ) ? ( n329 ) : ( n380 ) ;
assign n382 =  ( n322 ) ? ( n327 ) : ( n381 ) ;
assign n383 =  ( n320 ) ? ( n325 ) : ( n382 ) ;
assign n384 =  ( n332 ) ? ( n334 ) : ( n321 ) ;
assign n385 =  ( n330 ) ? ( n333 ) : ( n384 ) ;
assign n386 =  ( n328 ) ? ( n331 ) : ( n385 ) ;
assign n387 =  ( n326 ) ? ( n329 ) : ( n386 ) ;
assign n388 =  ( n324 ) ? ( n327 ) : ( n387 ) ;
assign n389 =  ( n322 ) ? ( n325 ) : ( n388 ) ;
assign n390 =  ( n320 ) ? ( n323 ) : ( n389 ) ;
assign n391 =  { ( n383 ) , ( n390 ) }  ;
assign n392 =  { ( n376 ) , ( n391 ) }  ;
assign n393 =  { ( n369 ) , ( n392 ) }  ;
assign n394 =  { ( n362 ) , ( n393 ) }  ;
assign n395 =  { ( n355 ) , ( n394 ) }  ;
assign n396 =  { ( n348 ) , ( n395 ) }  ;
assign n397 =  { ( n341 ) , ( n396 ) }  ;
assign n398 =  { ( n319 ) , ( n397 ) }  ;
assign n399 =  ( n42 ) ? ( slice_stream_buff_0 ) : ( n398 ) ;
assign n400 =  ( n9 ) ? ( slice_stream_buff_0 ) : ( slice_stream_buff_0 ) ;
assign n401 =  ( n44 ) ? ( n399 ) : ( n400 ) ;
assign n402 =  ( n37 ) ? ( slice_stream_buff_0 ) : ( n401 ) ;
assign n403 =  ( n30 ) ? ( slice_stream_buff_0 ) : ( n402 ) ;
assign n404 =  ( n4 ) ? ( slice_stream_buff_0 ) : ( n403 ) ;
assign n405 =  ( n21 ) ? ( slice_stream_buff_0 ) : ( n404 ) ;
assign n406 =  ( n42 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n407 =  ( n9 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_1 ) ;
assign n408 =  ( n44 ) ? ( n406 ) : ( n407 ) ;
assign n409 =  ( n37 ) ? ( slice_stream_buff_1 ) : ( n408 ) ;
assign n410 =  ( n30 ) ? ( slice_stream_buff_1 ) : ( n409 ) ;
assign n411 =  ( n4 ) ? ( slice_stream_buff_1 ) : ( n410 ) ;
assign n412 =  ( n21 ) ? ( slice_stream_buff_1 ) : ( n411 ) ;
assign n413 =  ( n86 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n414 =  ( n42 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n415 =  ( n9 ) ? ( slice_stream_empty ) : ( slice_stream_empty ) ;
assign n416 =  ( n44 ) ? ( n414 ) : ( n415 ) ;
assign n417 =  ( n37 ) ? ( n413 ) : ( n416 ) ;
assign n418 =  ( n30 ) ? ( slice_stream_empty ) : ( n417 ) ;
assign n419 =  ( n4 ) ? ( slice_stream_empty ) : ( n418 ) ;
assign n420 =  ( n21 ) ? ( slice_stream_empty ) : ( n419 ) ;
assign n421 =  ( slice_stream_empty ) == ( 1'd1 )  ;
assign n422 =  ( n421 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n423 =  ( n42 ) ? ( 1'd0 ) : ( n422 ) ;
assign n424 =  ( n9 ) ? ( slice_stream_full ) : ( slice_stream_full ) ;
assign n425 =  ( n44 ) ? ( n423 ) : ( n424 ) ;
assign n426 =  ( n37 ) ? ( 1'd0 ) : ( n425 ) ;
assign n427 =  ( n30 ) ? ( slice_stream_full ) : ( n426 ) ;
assign n428 =  ( n4 ) ? ( slice_stream_full ) : ( n427 ) ;
assign n429 =  ( n21 ) ? ( slice_stream_full ) : ( n428 ) ;
assign n430 =  ( LB2D_shift_x ) >= ( 9'd8 )  ;
assign n431 = n87[71:64] ;
assign n432 = LB2D_shift_0[71:64] ;
assign n433 = LB2D_shift_1[71:64] ;
assign n434 = LB2D_shift_2[71:64] ;
assign n435 = LB2D_shift_3[71:64] ;
assign n436 = LB2D_shift_4[71:64] ;
assign n437 = LB2D_shift_5[71:64] ;
assign n438 = LB2D_shift_6[71:64] ;
assign n439 = LB2D_shift_7[71:64] ;
assign n440 =  { ( n438 ) , ( n439 ) }  ;
assign n441 =  { ( n437 ) , ( n440 ) }  ;
assign n442 =  { ( n436 ) , ( n441 ) }  ;
assign n443 =  { ( n435 ) , ( n442 ) }  ;
assign n444 =  { ( n434 ) , ( n443 ) }  ;
assign n445 =  { ( n433 ) , ( n444 ) }  ;
assign n446 =  { ( n432 ) , ( n445 ) }  ;
assign n447 =  { ( n431 ) , ( n446 ) }  ;
assign n448 = n87[63:56] ;
assign n449 = LB2D_shift_0[63:56] ;
assign n450 = LB2D_shift_1[63:56] ;
assign n451 = LB2D_shift_2[63:56] ;
assign n452 = LB2D_shift_3[63:56] ;
assign n453 = LB2D_shift_4[63:56] ;
assign n454 = LB2D_shift_5[63:56] ;
assign n455 = LB2D_shift_6[63:56] ;
assign n456 = LB2D_shift_7[63:56] ;
assign n457 =  { ( n455 ) , ( n456 ) }  ;
assign n458 =  { ( n454 ) , ( n457 ) }  ;
assign n459 =  { ( n453 ) , ( n458 ) }  ;
assign n460 =  { ( n452 ) , ( n459 ) }  ;
assign n461 =  { ( n451 ) , ( n460 ) }  ;
assign n462 =  { ( n450 ) , ( n461 ) }  ;
assign n463 =  { ( n449 ) , ( n462 ) }  ;
assign n464 =  { ( n448 ) , ( n463 ) }  ;
assign n465 = n87[55:48] ;
assign n466 = LB2D_shift_0[55:48] ;
assign n467 = LB2D_shift_1[55:48] ;
assign n468 = LB2D_shift_2[55:48] ;
assign n469 = LB2D_shift_3[55:48] ;
assign n470 = LB2D_shift_4[55:48] ;
assign n471 = LB2D_shift_5[55:48] ;
assign n472 = LB2D_shift_6[55:48] ;
assign n473 = LB2D_shift_7[55:48] ;
assign n474 =  { ( n472 ) , ( n473 ) }  ;
assign n475 =  { ( n471 ) , ( n474 ) }  ;
assign n476 =  { ( n470 ) , ( n475 ) }  ;
assign n477 =  { ( n469 ) , ( n476 ) }  ;
assign n478 =  { ( n468 ) , ( n477 ) }  ;
assign n479 =  { ( n467 ) , ( n478 ) }  ;
assign n480 =  { ( n466 ) , ( n479 ) }  ;
assign n481 =  { ( n465 ) , ( n480 ) }  ;
assign n482 = n87[47:40] ;
assign n483 = LB2D_shift_0[47:40] ;
assign n484 = LB2D_shift_1[47:40] ;
assign n485 = LB2D_shift_2[47:40] ;
assign n486 = LB2D_shift_3[47:40] ;
assign n487 = LB2D_shift_4[47:40] ;
assign n488 = LB2D_shift_5[47:40] ;
assign n489 = LB2D_shift_6[47:40] ;
assign n490 = LB2D_shift_7[47:40] ;
assign n491 =  { ( n489 ) , ( n490 ) }  ;
assign n492 =  { ( n488 ) , ( n491 ) }  ;
assign n493 =  { ( n487 ) , ( n492 ) }  ;
assign n494 =  { ( n486 ) , ( n493 ) }  ;
assign n495 =  { ( n485 ) , ( n494 ) }  ;
assign n496 =  { ( n484 ) , ( n495 ) }  ;
assign n497 =  { ( n483 ) , ( n496 ) }  ;
assign n498 =  { ( n482 ) , ( n497 ) }  ;
assign n499 = n87[39:32] ;
assign n500 = LB2D_shift_0[39:32] ;
assign n501 = LB2D_shift_1[39:32] ;
assign n502 = LB2D_shift_2[39:32] ;
assign n503 = LB2D_shift_3[39:32] ;
assign n504 = LB2D_shift_4[39:32] ;
assign n505 = LB2D_shift_5[39:32] ;
assign n506 = LB2D_shift_6[39:32] ;
assign n507 = LB2D_shift_7[39:32] ;
assign n508 =  { ( n506 ) , ( n507 ) }  ;
assign n509 =  { ( n505 ) , ( n508 ) }  ;
assign n510 =  { ( n504 ) , ( n509 ) }  ;
assign n511 =  { ( n503 ) , ( n510 ) }  ;
assign n512 =  { ( n502 ) , ( n511 ) }  ;
assign n513 =  { ( n501 ) , ( n512 ) }  ;
assign n514 =  { ( n500 ) , ( n513 ) }  ;
assign n515 =  { ( n499 ) , ( n514 ) }  ;
assign n516 = n87[31:24] ;
assign n517 = LB2D_shift_0[31:24] ;
assign n518 = LB2D_shift_1[31:24] ;
assign n519 = LB2D_shift_2[31:24] ;
assign n520 = LB2D_shift_3[31:24] ;
assign n521 = LB2D_shift_4[31:24] ;
assign n522 = LB2D_shift_5[31:24] ;
assign n523 = LB2D_shift_6[31:24] ;
assign n524 = LB2D_shift_7[31:24] ;
assign n525 =  { ( n523 ) , ( n524 ) }  ;
assign n526 =  { ( n522 ) , ( n525 ) }  ;
assign n527 =  { ( n521 ) , ( n526 ) }  ;
assign n528 =  { ( n520 ) , ( n527 ) }  ;
assign n529 =  { ( n519 ) , ( n528 ) }  ;
assign n530 =  { ( n518 ) , ( n529 ) }  ;
assign n531 =  { ( n517 ) , ( n530 ) }  ;
assign n532 =  { ( n516 ) , ( n531 ) }  ;
assign n533 = n87[23:16] ;
assign n534 = LB2D_shift_0[23:16] ;
assign n535 = LB2D_shift_1[23:16] ;
assign n536 = LB2D_shift_2[23:16] ;
assign n537 = LB2D_shift_3[23:16] ;
assign n538 = LB2D_shift_4[23:16] ;
assign n539 = LB2D_shift_5[23:16] ;
assign n540 = LB2D_shift_6[23:16] ;
assign n541 = LB2D_shift_7[23:16] ;
assign n542 =  { ( n540 ) , ( n541 ) }  ;
assign n543 =  { ( n539 ) , ( n542 ) }  ;
assign n544 =  { ( n538 ) , ( n543 ) }  ;
assign n545 =  { ( n537 ) , ( n544 ) }  ;
assign n546 =  { ( n536 ) , ( n545 ) }  ;
assign n547 =  { ( n535 ) , ( n546 ) }  ;
assign n548 =  { ( n534 ) , ( n547 ) }  ;
assign n549 =  { ( n533 ) , ( n548 ) }  ;
assign n550 = n87[15:8] ;
assign n551 = LB2D_shift_0[15:8] ;
assign n552 = LB2D_shift_1[15:8] ;
assign n553 = LB2D_shift_2[15:8] ;
assign n554 = LB2D_shift_3[15:8] ;
assign n555 = LB2D_shift_4[15:8] ;
assign n556 = LB2D_shift_5[15:8] ;
assign n557 = LB2D_shift_6[15:8] ;
assign n558 = LB2D_shift_7[15:8] ;
assign n559 =  { ( n557 ) , ( n558 ) }  ;
assign n560 =  { ( n556 ) , ( n559 ) }  ;
assign n561 =  { ( n555 ) , ( n560 ) }  ;
assign n562 =  { ( n554 ) , ( n561 ) }  ;
assign n563 =  { ( n553 ) , ( n562 ) }  ;
assign n564 =  { ( n552 ) , ( n563 ) }  ;
assign n565 =  { ( n551 ) , ( n564 ) }  ;
assign n566 =  { ( n550 ) , ( n565 ) }  ;
assign n567 = n87[7:0] ;
assign n568 = LB2D_shift_0[7:0] ;
assign n569 = LB2D_shift_1[7:0] ;
assign n570 = LB2D_shift_2[7:0] ;
assign n571 = LB2D_shift_3[7:0] ;
assign n572 = LB2D_shift_4[7:0] ;
assign n573 = LB2D_shift_5[7:0] ;
assign n574 = LB2D_shift_6[7:0] ;
assign n575 = LB2D_shift_7[7:0] ;
assign n576 =  { ( n574 ) , ( n575 ) }  ;
assign n577 =  { ( n573 ) , ( n576 ) }  ;
assign n578 =  { ( n572 ) , ( n577 ) }  ;
assign n579 =  { ( n571 ) , ( n578 ) }  ;
assign n580 =  { ( n570 ) , ( n579 ) }  ;
assign n581 =  { ( n569 ) , ( n580 ) }  ;
assign n582 =  { ( n568 ) , ( n581 ) }  ;
assign n583 =  { ( n567 ) , ( n582 ) }  ;
assign n584 =  { ( n566 ) , ( n583 ) }  ;
assign n585 =  { ( n549 ) , ( n584 ) }  ;
assign n586 =  { ( n532 ) , ( n585 ) }  ;
assign n587 =  { ( n515 ) , ( n586 ) }  ;
assign n588 =  { ( n498 ) , ( n587 ) }  ;
assign n589 =  { ( n481 ) , ( n588 ) }  ;
assign n590 =  { ( n464 ) , ( n589 ) }  ;
assign n591 =  { ( n447 ) , ( n590 ) }  ;
assign n592 =  ( n430 ) ? ( n591 ) : ( stencil_stream_buff_0 ) ;
assign n593 =  ( n9 ) ? ( stencil_stream_buff_0 ) : ( stencil_stream_buff_0 ) ;
assign n594 =  ( n44 ) ? ( stencil_stream_buff_0 ) : ( n593 ) ;
assign n595 =  ( n37 ) ? ( n592 ) : ( n594 ) ;
assign n596 =  ( n30 ) ? ( stencil_stream_buff_0 ) : ( n595 ) ;
assign n597 =  ( n4 ) ? ( stencil_stream_buff_0 ) : ( n596 ) ;
assign n598 =  ( n21 ) ? ( stencil_stream_buff_0 ) : ( n597 ) ;
assign n599 =  ( n9 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_1 ) ;
assign n600 =  ( n44 ) ? ( stencil_stream_buff_1 ) : ( n599 ) ;
assign n601 =  ( n37 ) ? ( stencil_stream_buff_0 ) : ( n600 ) ;
assign n602 =  ( n30 ) ? ( stencil_stream_buff_1 ) : ( n601 ) ;
assign n603 =  ( n4 ) ? ( stencil_stream_buff_1 ) : ( n602 ) ;
assign n604 =  ( n21 ) ? ( stencil_stream_buff_1 ) : ( n603 ) ;
assign n605 =  ( n154 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n606 =  ( n35 ) ? ( stencil_stream_empty ) : ( 1'd0 ) ;
assign n607 =  ( n9 ) ? ( stencil_stream_empty ) : ( stencil_stream_empty ) ;
assign n608 =  ( n44 ) ? ( stencil_stream_empty ) : ( n607 ) ;
assign n609 =  ( n37 ) ? ( n606 ) : ( n608 ) ;
assign n610 =  ( n30 ) ? ( n605 ) : ( n609 ) ;
assign n611 =  ( n4 ) ? ( stencil_stream_empty ) : ( n610 ) ;
assign n612 =  ( n21 ) ? ( stencil_stream_empty ) : ( n611 ) ;
assign n613 =  ( n26 ) ? ( 1'd0 ) : ( 1'd0 ) ;
assign n614 =  ( stencil_stream_empty ) == ( 1'd1 )  ;
assign n615 =  ( n614 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n616 =  ( n35 ) ? ( stencil_stream_full ) : ( n615 ) ;
assign n617 =  ( n9 ) ? ( stencil_stream_full ) : ( stencil_stream_full ) ;
assign n618 =  ( n44 ) ? ( stencil_stream_full ) : ( n617 ) ;
assign n619 =  ( n37 ) ? ( n616 ) : ( n618 ) ;
assign n620 =  ( n30 ) ? ( n613 ) : ( n619 ) ;
assign n621 =  ( n4 ) ? ( stencil_stream_full ) : ( n620 ) ;
assign n622 =  ( n21 ) ? ( stencil_stream_full ) : ( n621 ) ;
assign n623 = ~ ( n21 ) ;
assign n624 = ~ ( n4 ) ;
assign n625 =  ( n623 ) & ( n624 )  ;
assign n626 = ~ ( n30 ) ;
assign n627 =  ( n625 ) & ( n626 )  ;
assign n628 = ~ ( n37 ) ;
assign n629 =  ( n627 ) & ( n628 )  ;
assign n630 = ~ ( n44 ) ;
assign n631 =  ( n629 ) & ( n630 )  ;
assign n632 = ~ ( n9 ) ;
assign n633 =  ( n631 ) & ( n632 )  ;
assign n634 =  ( n631 ) & ( n9 )  ;
assign n635 =  ( n629 ) & ( n44 )  ;
assign n636 = ~ ( n320 ) ;
assign n637 =  ( n635 ) & ( n636 )  ;
assign n638 =  ( n635 ) & ( n320 )  ;
assign n639 =  ( n627 ) & ( n37 )  ;
assign n640 =  ( n625 ) & ( n30 )  ;
assign n641 =  ( n623 ) & ( n4 )  ;
assign LB2D_proc_0_addr0 = n638 ? (LB2D_proc_x) : (0);
assign LB2D_proc_0_data0 = n638 ? (n319) : (LB2D_proc_0[0]);
assign n642 = ~ ( n322 ) ;
assign n643 =  ( n635 ) & ( n642 )  ;
assign n644 =  ( n635 ) & ( n322 )  ;
assign LB2D_proc_1_addr0 = n644 ? (LB2D_proc_x) : (0);
assign LB2D_proc_1_data0 = n644 ? (n319) : (LB2D_proc_1[0]);
assign n645 = ~ ( n324 ) ;
assign n646 =  ( n635 ) & ( n645 )  ;
assign n647 =  ( n635 ) & ( n324 )  ;
assign LB2D_proc_2_addr0 = n647 ? (LB2D_proc_x) : (0);
assign LB2D_proc_2_data0 = n647 ? (n319) : (LB2D_proc_2[0]);
assign n648 = ~ ( n326 ) ;
assign n649 =  ( n635 ) & ( n648 )  ;
assign n650 =  ( n635 ) & ( n326 )  ;
assign LB2D_proc_3_addr0 = n650 ? (LB2D_proc_x) : (0);
assign LB2D_proc_3_data0 = n650 ? (n319) : (LB2D_proc_3[0]);
assign n651 = ~ ( n328 ) ;
assign n652 =  ( n635 ) & ( n651 )  ;
assign n653 =  ( n635 ) & ( n328 )  ;
assign LB2D_proc_4_addr0 = n653 ? (LB2D_proc_x) : (0);
assign LB2D_proc_4_data0 = n653 ? (n319) : (LB2D_proc_4[0]);
assign n654 = ~ ( n330 ) ;
assign n655 =  ( n635 ) & ( n654 )  ;
assign n656 =  ( n635 ) & ( n330 )  ;
assign LB2D_proc_5_addr0 = n656 ? (LB2D_proc_x) : (0);
assign LB2D_proc_5_data0 = n656 ? (n319) : (LB2D_proc_5[0]);
assign n657 = ~ ( n332 ) ;
assign n658 =  ( n635 ) & ( n657 )  ;
assign n659 =  ( n635 ) & ( n332 )  ;
assign LB2D_proc_6_addr0 = n659 ? (LB2D_proc_x) : (0);
assign LB2D_proc_6_data0 = n659 ? (n319) : (LB2D_proc_6[0]);
assign n660 =  ( LB2D_proc_w ) == ( 64'd7 )  ;
assign n661 = ~ ( n660 ) ;
assign n662 =  ( n635 ) & ( n661 )  ;
assign n663 =  ( n635 ) & ( n660 )  ;
assign LB2D_proc_7_addr0 = n663 ? (LB2D_proc_x) : (0);
assign LB2D_proc_7_data0 = n663 ? (n319) : (LB2D_proc_7[0]);
/*
function [7:0] gb_fun ;
input [647:0] arg0;
    begin
//TODO: Add the specific function HERE.    end
endfunction
*/

always @(posedge clk) begin
   if(rst) begin
       LB1D_buff <= LB1D_buff;
       LB1D_in <= LB1D_in;
       LB1D_it_1 <= LB1D_it_1;
       LB1D_p_cnt <= LB1D_p_cnt;
       LB2D_proc_w <= LB2D_proc_w;
       LB2D_proc_x <= LB2D_proc_x;
       LB2D_proc_y <= LB2D_proc_y;
       LB2D_shift_0 <= LB2D_shift_0;
       LB2D_shift_1 <= LB2D_shift_1;
       LB2D_shift_2 <= LB2D_shift_2;
       LB2D_shift_3 <= LB2D_shift_3;
       LB2D_shift_4 <= LB2D_shift_4;
       LB2D_shift_5 <= LB2D_shift_5;
       LB2D_shift_6 <= LB2D_shift_6;
       LB2D_shift_7 <= LB2D_shift_7;
       LB2D_shift_x <= LB2D_shift_x;
       LB2D_shift_y <= LB2D_shift_y;
       arg_0_TDATA <= arg_0_TDATA;
       arg_0_TVALID <= arg_0_TVALID;
       arg_1_TREADY <= arg_1_TREADY;
       gb_exit_it_1 <= gb_exit_it_1;
       gb_exit_it_2 <= gb_exit_it_2;
       gb_exit_it_3 <= gb_exit_it_3;
       gb_exit_it_4 <= gb_exit_it_4;
       gb_exit_it_5 <= gb_exit_it_5;
       gb_exit_it_6 <= gb_exit_it_6;
       gb_exit_it_7 <= gb_exit_it_7;
       gb_exit_it_8 <= gb_exit_it_8;
       gb_p_cnt <= gb_p_cnt;
       gb_pp_it_1 <= gb_pp_it_1;
       gb_pp_it_2 <= gb_pp_it_2;
       gb_pp_it_3 <= gb_pp_it_3;
       gb_pp_it_4 <= gb_pp_it_4;
       gb_pp_it_5 <= gb_pp_it_5;
       gb_pp_it_6 <= gb_pp_it_6;
       gb_pp_it_7 <= gb_pp_it_7;
       gb_pp_it_8 <= gb_pp_it_8;
       gb_pp_it_9 <= gb_pp_it_9;
       in_stream_buff_0 <= in_stream_buff_0;
       in_stream_buff_1 <= in_stream_buff_1;
       in_stream_empty <= in_stream_empty;
       in_stream_full <= in_stream_full;
       slice_stream_buff_0 <= slice_stream_buff_0;
       slice_stream_buff_1 <= slice_stream_buff_1;
       slice_stream_empty <= slice_stream_empty;
       slice_stream_full <= slice_stream_full;
       stencil_stream_buff_0 <= stencil_stream_buff_0;
       stencil_stream_buff_1 <= stencil_stream_buff_1;
       stencil_stream_empty <= stencil_stream_empty;
       stencil_stream_full <= stencil_stream_full;
   end
   else if(step) begin
       LB1D_buff <= n11;
       LB1D_in <= n13;
       LB1D_it_1 <= n16;
       LB1D_p_cnt <= n55;
       LB2D_proc_w <= n66;
       LB2D_proc_x <= n77;
       LB2D_proc_y <= n85;
       LB2D_shift_0 <= n93;
       LB2D_shift_1 <= n99;
       LB2D_shift_2 <= n105;
       LB2D_shift_3 <= n111;
       LB2D_shift_4 <= n117;
       LB2D_shift_5 <= n123;
       LB2D_shift_6 <= n129;
       LB2D_shift_7 <= n135;
       LB2D_shift_x <= n142;
       LB2D_shift_y <= n153;
       arg_0_TDATA <= n162;
       arg_0_TVALID <= n170;
       arg_1_TREADY <= n177;
       gb_exit_it_1 <= n186;
       gb_exit_it_2 <= n192;
       gb_exit_it_3 <= n198;
       gb_exit_it_4 <= n204;
       gb_exit_it_5 <= n210;
       gb_exit_it_6 <= n216;
       gb_exit_it_7 <= n222;
       gb_exit_it_8 <= n228;
       gb_p_cnt <= n236;
       gb_pp_it_1 <= n242;
       gb_pp_it_2 <= n248;
       gb_pp_it_3 <= n254;
       gb_pp_it_4 <= n260;
       gb_pp_it_5 <= n266;
       gb_pp_it_6 <= n272;
       gb_pp_it_7 <= n278;
       gb_pp_it_8 <= n284;
       gb_pp_it_9 <= n290;
       in_stream_buff_0 <= n296;
       in_stream_buff_1 <= n302;
       in_stream_empty <= n310;
       in_stream_full <= n318;
       slice_stream_buff_0 <= n405;
       slice_stream_buff_1 <= n412;
       slice_stream_empty <= n420;
       slice_stream_full <= n429;
       stencil_stream_buff_0 <= n598;
       stencil_stream_buff_1 <= n604;
       stencil_stream_empty <= n612;
       stencil_stream_full <= n622;
       LB2D_proc_0 [ LB2D_proc_0_addr0 ] <= LB2D_proc_0_data0;
       LB2D_proc_1 [ LB2D_proc_1_addr0 ] <= LB2D_proc_1_data0;
       LB2D_proc_2 [ LB2D_proc_2_addr0 ] <= LB2D_proc_2_data0;
       LB2D_proc_3 [ LB2D_proc_3_addr0 ] <= LB2D_proc_3_data0;
       LB2D_proc_4 [ LB2D_proc_4_addr0 ] <= LB2D_proc_4_data0;
       LB2D_proc_5 [ LB2D_proc_5_addr0 ] <= LB2D_proc_5_data0;
       LB2D_proc_6 [ LB2D_proc_6_addr0 ] <= LB2D_proc_6_data0;
       LB2D_proc_7 [ LB2D_proc_7_addr0 ] <= LB2D_proc_7_data0;
   end
end
endmodule
