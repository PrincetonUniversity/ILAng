module gaussianRTL(
arg_0_TREADY,
arg_1_TDATA,
arg_1_TVALID,
LB2D_shift_0,
LB2D_shift_1,
LB2D_shift_2,
LB2D_shift_3,
LB2D_shift_4,
LB2D_shift_5,
LB2D_shift_6,
LB2D_shift_7,
LB2D_w_idx,
LB2D_x_idx,
LB2D_y_idx,
arg_0_TDATA,
arg_0_TVALID,
arg_1_TREADY,
slice_buff,
slice_full,
stencil_buff,
stencil_full,
clk,rst,
step
);
input            arg_0_TREADY;
input      [7:0] arg_1_TDATA;
input            arg_1_TVALID;
input clk;
input rst;
input step;
output     [71:0] LB2D_shift_0;
output     [71:0] LB2D_shift_1;
output     [71:0] LB2D_shift_2;
output     [71:0] LB2D_shift_3;
output     [71:0] LB2D_shift_4;
output     [71:0] LB2D_shift_5;
output     [71:0] LB2D_shift_6;
output     [71:0] LB2D_shift_7;
output     [63:0] LB2D_w_idx;
output      [8:0] LB2D_x_idx;
output      [9:0] LB2D_y_idx;
output      [7:0] arg_0_TDATA;
output            arg_0_TVALID;
output            arg_1_TREADY;
output     [71:0] slice_buff;
output            slice_full;
output    [647:0] stencil_buff;
output            stencil_full;
reg     [71:0] LB2D_shift_0;
reg     [71:0] LB2D_shift_1;
reg     [71:0] LB2D_shift_2;
reg     [71:0] LB2D_shift_3;
reg     [71:0] LB2D_shift_4;
reg     [71:0] LB2D_shift_5;
reg     [71:0] LB2D_shift_6;
reg     [71:0] LB2D_shift_7;
reg     [63:0] LB2D_w_idx;
reg      [8:0] LB2D_x_idx;
reg      [9:0] LB2D_y_idx;
reg      [7:0] arg_0_TDATA;
reg            arg_0_TVALID;
reg            arg_1_TREADY;
reg     [71:0] slice_buff;
reg            slice_full;
reg    [647:0] stencil_buff;
reg            stencil_full;
wire            arg_0_TREADY;
wire      [7:0] arg_1_TDATA;
wire            arg_1_TVALID;
wire            n0;
wire            n1;
wire            n2;
wire            n3;
wire            n4;
wire            n5;
wire            n6;
wire            n7;
wire            n8;
wire            n9;
wire            n10;
wire     [71:0] n11;
wire     [71:0] n12;
wire     [71:0] n13;
wire     [71:0] n14;
wire     [71:0] n15;
wire     [71:0] n16;
wire     [71:0] n17;
wire     [71:0] n18;
wire     [71:0] n19;
wire     [71:0] n20;
wire     [71:0] n21;
wire     [71:0] n22;
wire     [71:0] n23;
wire     [71:0] n24;
wire     [71:0] n25;
wire     [71:0] n26;
wire     [71:0] n27;
wire     [71:0] n28;
wire     [71:0] n29;
wire     [71:0] n30;
wire     [71:0] n31;
wire     [71:0] n32;
wire     [71:0] n33;
wire     [71:0] n34;
wire            n35;
wire            n36;
wire     [63:0] n37;
wire     [63:0] n38;
wire     [63:0] n39;
wire     [63:0] n40;
wire     [63:0] n41;
wire     [63:0] n42;
wire            n43;
wire      [8:0] n44;
wire      [8:0] n45;
wire      [8:0] n46;
wire      [8:0] n47;
wire      [8:0] n48;
wire            n49;
wire      [9:0] n50;
wire      [9:0] n51;
wire      [9:0] n52;
wire      [9:0] n53;
wire      [9:0] n54;
wire      [9:0] n55;
wire      [7:0] n56;
wire      [7:0] n57;
wire      [7:0] n58;
wire            n59;
wire            n60;
wire            n61;
wire            n62;
wire            n63;
wire            n64;
wire            n65;
wire            n66;
wire      [7:0] n67;
wire            n68;
wire      [7:0] n69;
wire            n70;
wire      [7:0] n71;
wire            n72;
wire      [7:0] n73;
wire            n74;
wire      [7:0] n75;
wire            n76;
wire      [7:0] n77;
wire            n78;
wire      [7:0] n79;
wire      [7:0] n80;
wire      [7:0] n81;
wire      [7:0] n82;
wire      [7:0] n83;
wire      [7:0] n84;
wire      [7:0] n85;
wire      [7:0] n86;
wire      [7:0] n87;
wire      [7:0] n88;
wire      [7:0] n89;
wire      [7:0] n90;
wire      [7:0] n91;
wire      [7:0] n92;
wire      [7:0] n93;
wire      [7:0] n94;
wire      [7:0] n95;
wire      [7:0] n96;
wire      [7:0] n97;
wire      [7:0] n98;
wire      [7:0] n99;
wire      [7:0] n100;
wire      [7:0] n101;
wire      [7:0] n102;
wire      [7:0] n103;
wire      [7:0] n104;
wire      [7:0] n105;
wire      [7:0] n106;
wire      [7:0] n107;
wire      [7:0] n108;
wire      [7:0] n109;
wire      [7:0] n110;
wire      [7:0] n111;
wire      [7:0] n112;
wire      [7:0] n113;
wire      [7:0] n114;
wire      [7:0] n115;
wire      [7:0] n116;
wire      [7:0] n117;
wire      [7:0] n118;
wire      [7:0] n119;
wire      [7:0] n120;
wire      [7:0] n121;
wire      [7:0] n122;
wire      [7:0] n123;
wire      [7:0] n124;
wire      [7:0] n125;
wire      [7:0] n126;
wire      [7:0] n127;
wire      [7:0] n128;
wire      [7:0] n129;
wire      [7:0] n130;
wire      [7:0] n131;
wire      [7:0] n132;
wire      [7:0] n133;
wire      [7:0] n134;
wire      [7:0] n135;
wire      [7:0] n136;
wire     [15:0] n137;
wire     [23:0] n138;
wire     [31:0] n139;
wire     [39:0] n140;
wire     [47:0] n141;
wire     [55:0] n142;
wire     [63:0] n143;
wire     [71:0] n144;
wire     [71:0] n145;
wire     [71:0] n146;
wire     [71:0] n147;
wire     [71:0] n148;
wire            n149;
wire            n150;
wire            n151;
wire      [7:0] n152;
wire      [7:0] n153;
wire      [7:0] n154;
wire      [7:0] n155;
wire      [7:0] n156;
wire      [7:0] n157;
wire      [7:0] n158;
wire      [7:0] n159;
wire      [7:0] n160;
wire     [15:0] n161;
wire     [23:0] n162;
wire     [31:0] n163;
wire     [39:0] n164;
wire     [47:0] n165;
wire     [55:0] n166;
wire     [63:0] n167;
wire     [71:0] n168;
wire      [7:0] n169;
wire      [7:0] n170;
wire      [7:0] n171;
wire      [7:0] n172;
wire      [7:0] n173;
wire      [7:0] n174;
wire      [7:0] n175;
wire      [7:0] n176;
wire      [7:0] n177;
wire     [15:0] n178;
wire     [23:0] n179;
wire     [31:0] n180;
wire     [39:0] n181;
wire     [47:0] n182;
wire     [55:0] n183;
wire     [63:0] n184;
wire     [71:0] n185;
wire      [7:0] n186;
wire      [7:0] n187;
wire      [7:0] n188;
wire      [7:0] n189;
wire      [7:0] n190;
wire      [7:0] n191;
wire      [7:0] n192;
wire      [7:0] n193;
wire      [7:0] n194;
wire     [15:0] n195;
wire     [23:0] n196;
wire     [31:0] n197;
wire     [39:0] n198;
wire     [47:0] n199;
wire     [55:0] n200;
wire     [63:0] n201;
wire     [71:0] n202;
wire      [7:0] n203;
wire      [7:0] n204;
wire      [7:0] n205;
wire      [7:0] n206;
wire      [7:0] n207;
wire      [7:0] n208;
wire      [7:0] n209;
wire      [7:0] n210;
wire      [7:0] n211;
wire     [15:0] n212;
wire     [23:0] n213;
wire     [31:0] n214;
wire     [39:0] n215;
wire     [47:0] n216;
wire     [55:0] n217;
wire     [63:0] n218;
wire     [71:0] n219;
wire      [7:0] n220;
wire      [7:0] n221;
wire      [7:0] n222;
wire      [7:0] n223;
wire      [7:0] n224;
wire      [7:0] n225;
wire      [7:0] n226;
wire      [7:0] n227;
wire      [7:0] n228;
wire     [15:0] n229;
wire     [23:0] n230;
wire     [31:0] n231;
wire     [39:0] n232;
wire     [47:0] n233;
wire     [55:0] n234;
wire     [63:0] n235;
wire     [71:0] n236;
wire      [7:0] n237;
wire      [7:0] n238;
wire      [7:0] n239;
wire      [7:0] n240;
wire      [7:0] n241;
wire      [7:0] n242;
wire      [7:0] n243;
wire      [7:0] n244;
wire      [7:0] n245;
wire     [15:0] n246;
wire     [23:0] n247;
wire     [31:0] n248;
wire     [39:0] n249;
wire     [47:0] n250;
wire     [55:0] n251;
wire     [63:0] n252;
wire     [71:0] n253;
wire      [7:0] n254;
wire      [7:0] n255;
wire      [7:0] n256;
wire      [7:0] n257;
wire      [7:0] n258;
wire      [7:0] n259;
wire      [7:0] n260;
wire      [7:0] n261;
wire      [7:0] n262;
wire     [15:0] n263;
wire     [23:0] n264;
wire     [31:0] n265;
wire     [39:0] n266;
wire     [47:0] n267;
wire     [55:0] n268;
wire     [63:0] n269;
wire     [71:0] n270;
wire      [7:0] n271;
wire      [7:0] n272;
wire      [7:0] n273;
wire      [7:0] n274;
wire      [7:0] n275;
wire      [7:0] n276;
wire      [7:0] n277;
wire      [7:0] n278;
wire      [7:0] n279;
wire     [15:0] n280;
wire     [23:0] n281;
wire     [31:0] n282;
wire     [39:0] n283;
wire     [47:0] n284;
wire     [55:0] n285;
wire     [63:0] n286;
wire     [71:0] n287;
wire      [7:0] n288;
wire      [7:0] n289;
wire      [7:0] n290;
wire      [7:0] n291;
wire      [7:0] n292;
wire      [7:0] n293;
wire      [7:0] n294;
wire      [7:0] n295;
wire      [7:0] n296;
wire     [15:0] n297;
wire     [23:0] n298;
wire     [31:0] n299;
wire     [39:0] n300;
wire     [47:0] n301;
wire     [55:0] n302;
wire     [63:0] n303;
wire     [71:0] n304;
wire    [143:0] n305;
wire    [215:0] n306;
wire    [287:0] n307;
wire    [359:0] n308;
wire    [431:0] n309;
wire    [503:0] n310;
wire    [575:0] n311;
wire    [647:0] n312;
wire    [647:0] n313;
wire    [647:0] n314;
wire    [647:0] n315;
wire            n316;
wire            n317;
wire            n318;
wire      [8:0] LB2D_buff_0_addr0;
wire      [7:0] LB2D_buff_0_data0;
wire            n319;
wire            n320;
wire            n321;
wire            n322;
wire            n323;
wire            n324;
wire            n325;
wire            n326;
wire            n327;
wire            n328;
wire      [8:0] LB2D_buff_1_addr0;
wire      [7:0] LB2D_buff_1_data0;
wire            n329;
wire            n330;
wire            n331;
wire      [8:0] LB2D_buff_2_addr0;
wire      [7:0] LB2D_buff_2_data0;
wire            n332;
wire            n333;
wire            n334;
wire      [8:0] LB2D_buff_3_addr0;
wire      [7:0] LB2D_buff_3_data0;
wire            n335;
wire            n336;
wire            n337;
wire      [8:0] LB2D_buff_4_addr0;
wire      [7:0] LB2D_buff_4_data0;
wire            n338;
wire            n339;
wire            n340;
wire      [8:0] LB2D_buff_5_addr0;
wire      [7:0] LB2D_buff_5_data0;
wire            n341;
wire            n342;
wire            n343;
wire      [8:0] LB2D_buff_6_addr0;
wire      [7:0] LB2D_buff_6_data0;
wire            n344;
wire            n345;
wire            n346;
wire      [8:0] LB2D_buff_7_addr0;
wire      [7:0] LB2D_buff_7_data0;
wire            n347;
wire            n348;
wire            n349;
wire            n350;
reg      [7:0] LB2D_buff_0[511:0];
reg      [7:0] LB2D_buff_1[511:0];
reg      [7:0] LB2D_buff_2[511:0];
reg      [7:0] LB2D_buff_3[511:0];
reg      [7:0] LB2D_buff_4[511:0];
reg      [7:0] LB2D_buff_5[511:0];
reg      [7:0] LB2D_buff_6[511:0];
reg      [7:0] LB2D_buff_7[511:0];
wire clk;
wire rst;
wire step;
assign n0 =  ( arg_1_TVALID ) == ( 1'd1 )  ;
assign n1 =  ( slice_full ) == ( 1'd0 )  ;
assign n2 =  ( n0 ) & ( n1 )  ;
assign n3 =  ( slice_full ) == ( 1'd1 )  ;
assign n4 =  ( stencil_full ) == ( 1'd0 )  ;
assign n5 =  ( n3 ) & ( n4 )  ;
assign n6 =  ( arg_0_TREADY ) == ( 1'd1 )  ;
assign n7 =  ( arg_0_TVALID ) == ( 1'd1 )  ;
assign n8 =  ( n6 ) & ( n7 )  ;
assign n9 =  ( arg_1_TVALID ) == ( 1'd0 )  ;
assign n10 =  ( n8 ) & ( n9 )  ;
assign n11 =  ( n10 ) ? ( LB2D_shift_0 ) : ( LB2D_shift_0 ) ;
assign n12 =  ( n5 ) ? ( slice_buff ) : ( n11 ) ;
assign n13 =  ( n2 ) ? ( LB2D_shift_0 ) : ( n12 ) ;
assign n14 =  ( n10 ) ? ( LB2D_shift_1 ) : ( LB2D_shift_1 ) ;
assign n15 =  ( n5 ) ? ( LB2D_shift_0 ) : ( n14 ) ;
assign n16 =  ( n2 ) ? ( LB2D_shift_1 ) : ( n15 ) ;
assign n17 =  ( n10 ) ? ( LB2D_shift_2 ) : ( LB2D_shift_2 ) ;
assign n18 =  ( n5 ) ? ( LB2D_shift_1 ) : ( n17 ) ;
assign n19 =  ( n2 ) ? ( LB2D_shift_2 ) : ( n18 ) ;
assign n20 =  ( n10 ) ? ( LB2D_shift_3 ) : ( LB2D_shift_3 ) ;
assign n21 =  ( n5 ) ? ( LB2D_shift_2 ) : ( n20 ) ;
assign n22 =  ( n2 ) ? ( LB2D_shift_3 ) : ( n21 ) ;
assign n23 =  ( n10 ) ? ( LB2D_shift_4 ) : ( LB2D_shift_4 ) ;
assign n24 =  ( n5 ) ? ( LB2D_shift_3 ) : ( n23 ) ;
assign n25 =  ( n2 ) ? ( LB2D_shift_4 ) : ( n24 ) ;
assign n26 =  ( n10 ) ? ( LB2D_shift_5 ) : ( LB2D_shift_5 ) ;
assign n27 =  ( n5 ) ? ( LB2D_shift_4 ) : ( n26 ) ;
assign n28 =  ( n2 ) ? ( LB2D_shift_5 ) : ( n27 ) ;
assign n29 =  ( n10 ) ? ( LB2D_shift_6 ) : ( LB2D_shift_6 ) ;
assign n30 =  ( n5 ) ? ( LB2D_shift_5 ) : ( n29 ) ;
assign n31 =  ( n2 ) ? ( LB2D_shift_6 ) : ( n30 ) ;
assign n32 =  ( n10 ) ? ( LB2D_shift_7 ) : ( LB2D_shift_7 ) ;
assign n33 =  ( n5 ) ? ( LB2D_shift_6 ) : ( n32 ) ;
assign n34 =  ( n2 ) ? ( LB2D_shift_7 ) : ( n33 ) ;
assign n35 =  ( LB2D_x_idx ) == ( 9'd487 )  ;
assign n36 =  ( LB2D_w_idx ) != ( 64'd7 )  ;
assign n37 =  ( LB2D_w_idx ) + ( 64'd1 )  ;
assign n38 =  ( n36 ) ? ( n37 ) : ( 64'd0 ) ;
assign n39 =  ( n35 ) ? ( n38 ) : ( LB2D_w_idx ) ;
assign n40 =  ( n10 ) ? ( LB2D_w_idx ) : ( LB2D_w_idx ) ;
assign n41 =  ( n5 ) ? ( LB2D_w_idx ) : ( n40 ) ;
assign n42 =  ( n2 ) ? ( n39 ) : ( n41 ) ;
assign n43 =  ( LB2D_x_idx ) != ( 9'd487 )  ;
assign n44 =  ( LB2D_x_idx ) + ( 9'd1 )  ;
assign n45 =  ( n43 ) ? ( n44 ) : ( 9'd0 ) ;
assign n46 =  ( n10 ) ? ( LB2D_x_idx ) : ( LB2D_x_idx ) ;
assign n47 =  ( n5 ) ? ( LB2D_x_idx ) : ( n46 ) ;
assign n48 =  ( n2 ) ? ( n45 ) : ( n47 ) ;
assign n49 =  ( LB2D_y_idx ) != ( 10'd687 )  ;
assign n50 =  ( LB2D_y_idx ) + ( 10'd1 )  ;
assign n51 =  ( n49 ) ? ( n50 ) : ( LB2D_y_idx ) ;
assign n52 =  ( n35 ) ? ( n51 ) : ( LB2D_y_idx ) ;
assign n53 =  ( n10 ) ? ( LB2D_y_idx ) : ( LB2D_y_idx ) ;
assign n54 =  ( n5 ) ? ( LB2D_y_idx ) : ( n53 ) ;
assign n55 =  ( n2 ) ? ( n52 ) : ( n54 ) ;
assign n56 =  ( n10 ) ? ( arg_0_TDATA ) : ( arg_0_TDATA ) ;
assign n57 =  ( n5 ) ? ( arg_0_TDATA ) : ( n56 ) ;
assign n58 =  ( n2 ) ? ( arg_0_TDATA ) : ( n57 ) ;
assign n59 =  ( n10 ) ? ( 1'd0 ) : ( arg_0_TVALID ) ;
assign n60 =  ( n5 ) ? ( 1'd0 ) : ( n59 ) ;
assign n61 =  ( n2 ) ? ( 1'd0 ) : ( n60 ) ;
assign n62 =  ( n10 ) ? ( 1'd1 ) : ( arg_1_TREADY ) ;
assign n63 =  ( n5 ) ? ( 1'd1 ) : ( n62 ) ;
assign n64 =  ( n2 ) ? ( 1'd0 ) : ( n63 ) ;
assign n65 =  ( LB2D_y_idx ) >= ( 10'd8 )  ;
assign n66 =  ( LB2D_w_idx ) == ( 64'd0 )  ;
assign n67 =  (  LB2D_buff_7 [ LB2D_x_idx ] )  ;
assign n68 =  ( LB2D_w_idx ) == ( 64'd1 )  ;
assign n69 =  (  LB2D_buff_0 [ LB2D_x_idx ] )  ;
assign n70 =  ( LB2D_w_idx ) == ( 64'd2 )  ;
assign n71 =  (  LB2D_buff_1 [ LB2D_x_idx ] )  ;
assign n72 =  ( LB2D_w_idx ) == ( 64'd3 )  ;
assign n73 =  (  LB2D_buff_2 [ LB2D_x_idx ] )  ;
assign n74 =  ( LB2D_w_idx ) == ( 64'd4 )  ;
assign n75 =  (  LB2D_buff_3 [ LB2D_x_idx ] )  ;
assign n76 =  ( LB2D_w_idx ) == ( 64'd5 )  ;
assign n77 =  (  LB2D_buff_4 [ LB2D_x_idx ] )  ;
assign n78 =  ( LB2D_w_idx ) == ( 64'd6 )  ;
assign n79 =  (  LB2D_buff_5 [ LB2D_x_idx ] )  ;
assign n80 =  (  LB2D_buff_6 [ LB2D_x_idx ] )  ;
assign n81 =  ( n78 ) ? ( n79 ) : ( n80 ) ;
assign n82 =  ( n76 ) ? ( n77 ) : ( n81 ) ;
assign n83 =  ( n74 ) ? ( n75 ) : ( n82 ) ;
assign n84 =  ( n72 ) ? ( n73 ) : ( n83 ) ;
assign n85 =  ( n70 ) ? ( n71 ) : ( n84 ) ;
assign n86 =  ( n68 ) ? ( n69 ) : ( n85 ) ;
assign n87 =  ( n66 ) ? ( n67 ) : ( n86 ) ;
assign n88 =  ( n78 ) ? ( n77 ) : ( n79 ) ;
assign n89 =  ( n76 ) ? ( n75 ) : ( n88 ) ;
assign n90 =  ( n74 ) ? ( n73 ) : ( n89 ) ;
assign n91 =  ( n72 ) ? ( n71 ) : ( n90 ) ;
assign n92 =  ( n70 ) ? ( n69 ) : ( n91 ) ;
assign n93 =  ( n68 ) ? ( n67 ) : ( n92 ) ;
assign n94 =  ( n66 ) ? ( n80 ) : ( n93 ) ;
assign n95 =  ( n78 ) ? ( n75 ) : ( n77 ) ;
assign n96 =  ( n76 ) ? ( n73 ) : ( n95 ) ;
assign n97 =  ( n74 ) ? ( n71 ) : ( n96 ) ;
assign n98 =  ( n72 ) ? ( n69 ) : ( n97 ) ;
assign n99 =  ( n70 ) ? ( n67 ) : ( n98 ) ;
assign n100 =  ( n68 ) ? ( n80 ) : ( n99 ) ;
assign n101 =  ( n66 ) ? ( n79 ) : ( n100 ) ;
assign n102 =  ( n78 ) ? ( n73 ) : ( n75 ) ;
assign n103 =  ( n76 ) ? ( n71 ) : ( n102 ) ;
assign n104 =  ( n74 ) ? ( n69 ) : ( n103 ) ;
assign n105 =  ( n72 ) ? ( n67 ) : ( n104 ) ;
assign n106 =  ( n70 ) ? ( n80 ) : ( n105 ) ;
assign n107 =  ( n68 ) ? ( n79 ) : ( n106 ) ;
assign n108 =  ( n66 ) ? ( n77 ) : ( n107 ) ;
assign n109 =  ( n78 ) ? ( n71 ) : ( n73 ) ;
assign n110 =  ( n76 ) ? ( n69 ) : ( n109 ) ;
assign n111 =  ( n74 ) ? ( n67 ) : ( n110 ) ;
assign n112 =  ( n72 ) ? ( n80 ) : ( n111 ) ;
assign n113 =  ( n70 ) ? ( n79 ) : ( n112 ) ;
assign n114 =  ( n68 ) ? ( n77 ) : ( n113 ) ;
assign n115 =  ( n66 ) ? ( n75 ) : ( n114 ) ;
assign n116 =  ( n78 ) ? ( n69 ) : ( n71 ) ;
assign n117 =  ( n76 ) ? ( n67 ) : ( n116 ) ;
assign n118 =  ( n74 ) ? ( n80 ) : ( n117 ) ;
assign n119 =  ( n72 ) ? ( n79 ) : ( n118 ) ;
assign n120 =  ( n70 ) ? ( n77 ) : ( n119 ) ;
assign n121 =  ( n68 ) ? ( n75 ) : ( n120 ) ;
assign n122 =  ( n66 ) ? ( n73 ) : ( n121 ) ;
assign n123 =  ( n78 ) ? ( n67 ) : ( n69 ) ;
assign n124 =  ( n76 ) ? ( n80 ) : ( n123 ) ;
assign n125 =  ( n74 ) ? ( n79 ) : ( n124 ) ;
assign n126 =  ( n72 ) ? ( n77 ) : ( n125 ) ;
assign n127 =  ( n70 ) ? ( n75 ) : ( n126 ) ;
assign n128 =  ( n68 ) ? ( n73 ) : ( n127 ) ;
assign n129 =  ( n66 ) ? ( n71 ) : ( n128 ) ;
assign n130 =  ( n78 ) ? ( n80 ) : ( n67 ) ;
assign n131 =  ( n76 ) ? ( n79 ) : ( n130 ) ;
assign n132 =  ( n74 ) ? ( n77 ) : ( n131 ) ;
assign n133 =  ( n72 ) ? ( n75 ) : ( n132 ) ;
assign n134 =  ( n70 ) ? ( n73 ) : ( n133 ) ;
assign n135 =  ( n68 ) ? ( n71 ) : ( n134 ) ;
assign n136 =  ( n66 ) ? ( n69 ) : ( n135 ) ;
assign n137 =  { ( n129 ) , ( n136 ) }  ;
assign n138 =  { ( n122 ) , ( n137 ) }  ;
assign n139 =  { ( n115 ) , ( n138 ) }  ;
assign n140 =  { ( n108 ) , ( n139 ) }  ;
assign n141 =  { ( n101 ) , ( n140 ) }  ;
assign n142 =  { ( n94 ) , ( n141 ) }  ;
assign n143 =  { ( n87 ) , ( n142 ) }  ;
assign n144 =  { ( arg_1_TDATA ) , ( n143 ) }  ;
assign n145 =  ( n65 ) ? ( n144 ) : ( slice_buff ) ;
assign n146 =  ( n10 ) ? ( slice_buff ) : ( slice_buff ) ;
assign n147 =  ( n5 ) ? ( slice_buff ) : ( n146 ) ;
assign n148 =  ( n2 ) ? ( n145 ) : ( n147 ) ;
assign n149 =  ( n10 ) ? ( slice_full ) : ( slice_full ) ;
assign n150 =  ( n5 ) ? ( 1'd0 ) : ( n149 ) ;
assign n151 =  ( n2 ) ? ( 1'd1 ) : ( n150 ) ;
assign n152 = slice_buff[71:64] ;
assign n153 = LB2D_shift_0[71:64] ;
assign n154 = LB2D_shift_1[71:64] ;
assign n155 = LB2D_shift_2[71:64] ;
assign n156 = LB2D_shift_3[71:64] ;
assign n157 = LB2D_shift_4[71:64] ;
assign n158 = LB2D_shift_5[71:64] ;
assign n159 = LB2D_shift_6[71:64] ;
assign n160 = LB2D_shift_7[71:64] ;
assign n161 =  { ( n159 ) , ( n160 ) }  ;
assign n162 =  { ( n158 ) , ( n161 ) }  ;
assign n163 =  { ( n157 ) , ( n162 ) }  ;
assign n164 =  { ( n156 ) , ( n163 ) }  ;
assign n165 =  { ( n155 ) , ( n164 ) }  ;
assign n166 =  { ( n154 ) , ( n165 ) }  ;
assign n167 =  { ( n153 ) , ( n166 ) }  ;
assign n168 =  { ( n152 ) , ( n167 ) }  ;
assign n169 = slice_buff[63:56] ;
assign n170 = LB2D_shift_0[63:56] ;
assign n171 = LB2D_shift_1[63:56] ;
assign n172 = LB2D_shift_2[63:56] ;
assign n173 = LB2D_shift_3[63:56] ;
assign n174 = LB2D_shift_4[63:56] ;
assign n175 = LB2D_shift_5[63:56] ;
assign n176 = LB2D_shift_6[63:56] ;
assign n177 = LB2D_shift_7[63:56] ;
assign n178 =  { ( n176 ) , ( n177 ) }  ;
assign n179 =  { ( n175 ) , ( n178 ) }  ;
assign n180 =  { ( n174 ) , ( n179 ) }  ;
assign n181 =  { ( n173 ) , ( n180 ) }  ;
assign n182 =  { ( n172 ) , ( n181 ) }  ;
assign n183 =  { ( n171 ) , ( n182 ) }  ;
assign n184 =  { ( n170 ) , ( n183 ) }  ;
assign n185 =  { ( n169 ) , ( n184 ) }  ;
assign n186 = slice_buff[55:48] ;
assign n187 = LB2D_shift_0[55:48] ;
assign n188 = LB2D_shift_1[55:48] ;
assign n189 = LB2D_shift_2[55:48] ;
assign n190 = LB2D_shift_3[55:48] ;
assign n191 = LB2D_shift_4[55:48] ;
assign n192 = LB2D_shift_5[55:48] ;
assign n193 = LB2D_shift_6[55:48] ;
assign n194 = LB2D_shift_7[55:48] ;
assign n195 =  { ( n193 ) , ( n194 ) }  ;
assign n196 =  { ( n192 ) , ( n195 ) }  ;
assign n197 =  { ( n191 ) , ( n196 ) }  ;
assign n198 =  { ( n190 ) , ( n197 ) }  ;
assign n199 =  { ( n189 ) , ( n198 ) }  ;
assign n200 =  { ( n188 ) , ( n199 ) }  ;
assign n201 =  { ( n187 ) , ( n200 ) }  ;
assign n202 =  { ( n186 ) , ( n201 ) }  ;
assign n203 = slice_buff[47:40] ;
assign n204 = LB2D_shift_0[47:40] ;
assign n205 = LB2D_shift_1[47:40] ;
assign n206 = LB2D_shift_2[47:40] ;
assign n207 = LB2D_shift_3[47:40] ;
assign n208 = LB2D_shift_4[47:40] ;
assign n209 = LB2D_shift_5[47:40] ;
assign n210 = LB2D_shift_6[47:40] ;
assign n211 = LB2D_shift_7[47:40] ;
assign n212 =  { ( n210 ) , ( n211 ) }  ;
assign n213 =  { ( n209 ) , ( n212 ) }  ;
assign n214 =  { ( n208 ) , ( n213 ) }  ;
assign n215 =  { ( n207 ) , ( n214 ) }  ;
assign n216 =  { ( n206 ) , ( n215 ) }  ;
assign n217 =  { ( n205 ) , ( n216 ) }  ;
assign n218 =  { ( n204 ) , ( n217 ) }  ;
assign n219 =  { ( n203 ) , ( n218 ) }  ;
assign n220 = slice_buff[39:32] ;
assign n221 = LB2D_shift_0[39:32] ;
assign n222 = LB2D_shift_1[39:32] ;
assign n223 = LB2D_shift_2[39:32] ;
assign n224 = LB2D_shift_3[39:32] ;
assign n225 = LB2D_shift_4[39:32] ;
assign n226 = LB2D_shift_5[39:32] ;
assign n227 = LB2D_shift_6[39:32] ;
assign n228 = LB2D_shift_7[39:32] ;
assign n229 =  { ( n227 ) , ( n228 ) }  ;
assign n230 =  { ( n226 ) , ( n229 ) }  ;
assign n231 =  { ( n225 ) , ( n230 ) }  ;
assign n232 =  { ( n224 ) , ( n231 ) }  ;
assign n233 =  { ( n223 ) , ( n232 ) }  ;
assign n234 =  { ( n222 ) , ( n233 ) }  ;
assign n235 =  { ( n221 ) , ( n234 ) }  ;
assign n236 =  { ( n220 ) , ( n235 ) }  ;
assign n237 = slice_buff[31:24] ;
assign n238 = LB2D_shift_0[31:24] ;
assign n239 = LB2D_shift_1[31:24] ;
assign n240 = LB2D_shift_2[31:24] ;
assign n241 = LB2D_shift_3[31:24] ;
assign n242 = LB2D_shift_4[31:24] ;
assign n243 = LB2D_shift_5[31:24] ;
assign n244 = LB2D_shift_6[31:24] ;
assign n245 = LB2D_shift_7[31:24] ;
assign n246 =  { ( n244 ) , ( n245 ) }  ;
assign n247 =  { ( n243 ) , ( n246 ) }  ;
assign n248 =  { ( n242 ) , ( n247 ) }  ;
assign n249 =  { ( n241 ) , ( n248 ) }  ;
assign n250 =  { ( n240 ) , ( n249 ) }  ;
assign n251 =  { ( n239 ) , ( n250 ) }  ;
assign n252 =  { ( n238 ) , ( n251 ) }  ;
assign n253 =  { ( n237 ) , ( n252 ) }  ;
assign n254 = slice_buff[23:16] ;
assign n255 = LB2D_shift_0[23:16] ;
assign n256 = LB2D_shift_1[23:16] ;
assign n257 = LB2D_shift_2[23:16] ;
assign n258 = LB2D_shift_3[23:16] ;
assign n259 = LB2D_shift_4[23:16] ;
assign n260 = LB2D_shift_5[23:16] ;
assign n261 = LB2D_shift_6[23:16] ;
assign n262 = LB2D_shift_7[23:16] ;
assign n263 =  { ( n261 ) , ( n262 ) }  ;
assign n264 =  { ( n260 ) , ( n263 ) }  ;
assign n265 =  { ( n259 ) , ( n264 ) }  ;
assign n266 =  { ( n258 ) , ( n265 ) }  ;
assign n267 =  { ( n257 ) , ( n266 ) }  ;
assign n268 =  { ( n256 ) , ( n267 ) }  ;
assign n269 =  { ( n255 ) , ( n268 ) }  ;
assign n270 =  { ( n254 ) , ( n269 ) }  ;
assign n271 = slice_buff[15:8] ;
assign n272 = LB2D_shift_0[15:8] ;
assign n273 = LB2D_shift_1[15:8] ;
assign n274 = LB2D_shift_2[15:8] ;
assign n275 = LB2D_shift_3[15:8] ;
assign n276 = LB2D_shift_4[15:8] ;
assign n277 = LB2D_shift_5[15:8] ;
assign n278 = LB2D_shift_6[15:8] ;
assign n279 = LB2D_shift_7[15:8] ;
assign n280 =  { ( n278 ) , ( n279 ) }  ;
assign n281 =  { ( n277 ) , ( n280 ) }  ;
assign n282 =  { ( n276 ) , ( n281 ) }  ;
assign n283 =  { ( n275 ) , ( n282 ) }  ;
assign n284 =  { ( n274 ) , ( n283 ) }  ;
assign n285 =  { ( n273 ) , ( n284 ) }  ;
assign n286 =  { ( n272 ) , ( n285 ) }  ;
assign n287 =  { ( n271 ) , ( n286 ) }  ;
assign n288 = slice_buff[7:0] ;
assign n289 = LB2D_shift_0[7:0] ;
assign n290 = LB2D_shift_1[7:0] ;
assign n291 = LB2D_shift_2[7:0] ;
assign n292 = LB2D_shift_3[7:0] ;
assign n293 = LB2D_shift_4[7:0] ;
assign n294 = LB2D_shift_5[7:0] ;
assign n295 = LB2D_shift_6[7:0] ;
assign n296 = LB2D_shift_7[7:0] ;
assign n297 =  { ( n295 ) , ( n296 ) }  ;
assign n298 =  { ( n294 ) , ( n297 ) }  ;
assign n299 =  { ( n293 ) , ( n298 ) }  ;
assign n300 =  { ( n292 ) , ( n299 ) }  ;
assign n301 =  { ( n291 ) , ( n300 ) }  ;
assign n302 =  { ( n290 ) , ( n301 ) }  ;
assign n303 =  { ( n289 ) , ( n302 ) }  ;
assign n304 =  { ( n288 ) , ( n303 ) }  ;
assign n305 =  { ( n287 ) , ( n304 ) }  ;
assign n306 =  { ( n270 ) , ( n305 ) }  ;
assign n307 =  { ( n253 ) , ( n306 ) }  ;
assign n308 =  { ( n236 ) , ( n307 ) }  ;
assign n309 =  { ( n219 ) , ( n308 ) }  ;
assign n310 =  { ( n202 ) , ( n309 ) }  ;
assign n311 =  { ( n185 ) , ( n310 ) }  ;
assign n312 =  { ( n168 ) , ( n311 ) }  ;
assign n313 =  ( n10 ) ? ( stencil_buff ) : ( stencil_buff ) ;
assign n314 =  ( n5 ) ? ( n312 ) : ( n313 ) ;
assign n315 =  ( n2 ) ? ( stencil_buff ) : ( n314 ) ;
assign n316 =  ( n10 ) ? ( 1'd0 ) : ( stencil_full ) ;
assign n317 =  ( n5 ) ? ( 1'd0 ) : ( n316 ) ;
assign n318 =  ( n2 ) ? ( stencil_full ) : ( n317 ) ;
assign n319 = ~ ( n2 ) ;
assign n320 = ~ ( n5 ) ;
assign n321 =  ( n319 ) & ( n320 )  ;
assign n322 = ~ ( n10 ) ;
assign n323 =  ( n321 ) & ( n322 )  ;
assign n324 =  ( n321 ) & ( n10 )  ;
assign n325 =  ( n319 ) & ( n5 )  ;
assign n326 = ~ ( n66 ) ;
assign n327 =  ( n2 ) & ( n326 )  ;
assign n328 =  ( n2 ) & ( n66 )  ;
assign LB2D_buff_0_addr0 = n328 ? (LB2D_x_idx) : (0);
assign LB2D_buff_0_data0 = n328 ? (arg_1_TDATA) : (LB2D_buff_0[0]);
assign n329 = ~ ( n68 ) ;
assign n330 =  ( n2 ) & ( n329 )  ;
assign n331 =  ( n2 ) & ( n68 )  ;
assign LB2D_buff_1_addr0 = n331 ? (LB2D_x_idx) : (0);
assign LB2D_buff_1_data0 = n331 ? (arg_1_TDATA) : (LB2D_buff_1[0]);
assign n332 = ~ ( n70 ) ;
assign n333 =  ( n2 ) & ( n332 )  ;
assign n334 =  ( n2 ) & ( n70 )  ;
assign LB2D_buff_2_addr0 = n334 ? (LB2D_x_idx) : (0);
assign LB2D_buff_2_data0 = n334 ? (arg_1_TDATA) : (LB2D_buff_2[0]);
assign n335 = ~ ( n72 ) ;
assign n336 =  ( n2 ) & ( n335 )  ;
assign n337 =  ( n2 ) & ( n72 )  ;
assign LB2D_buff_3_addr0 = n337 ? (LB2D_x_idx) : (0);
assign LB2D_buff_3_data0 = n337 ? (arg_1_TDATA) : (LB2D_buff_3[0]);
assign n338 = ~ ( n74 ) ;
assign n339 =  ( n2 ) & ( n338 )  ;
assign n340 =  ( n2 ) & ( n74 )  ;
assign LB2D_buff_4_addr0 = n340 ? (LB2D_x_idx) : (0);
assign LB2D_buff_4_data0 = n340 ? (arg_1_TDATA) : (LB2D_buff_4[0]);
assign n341 = ~ ( n76 ) ;
assign n342 =  ( n2 ) & ( n341 )  ;
assign n343 =  ( n2 ) & ( n76 )  ;
assign LB2D_buff_5_addr0 = n343 ? (LB2D_x_idx) : (0);
assign LB2D_buff_5_data0 = n343 ? (arg_1_TDATA) : (LB2D_buff_5[0]);
assign n344 = ~ ( n78 ) ;
assign n345 =  ( n2 ) & ( n344 )  ;
assign n346 =  ( n2 ) & ( n78 )  ;
assign LB2D_buff_6_addr0 = n346 ? (LB2D_x_idx) : (0);
assign LB2D_buff_6_data0 = n346 ? (arg_1_TDATA) : (LB2D_buff_6[0]);
assign n347 =  ( LB2D_w_idx ) == ( 64'd7 )  ;
assign n348 = ~ ( n347 ) ;
assign n349 =  ( n2 ) & ( n348 )  ;
assign n350 =  ( n2 ) & ( n347 )  ;
assign LB2D_buff_7_addr0 = n350 ? (LB2D_x_idx) : (0);
assign LB2D_buff_7_data0 = n350 ? (arg_1_TDATA) : (LB2D_buff_7[0]);
function [7:0] gaussianBlurStencil ;
input [647:0] arg0;
    begin
//TODO: Add the specific function HERE.    end
endfunction

always @(posedge clk) begin
   if(rst) begin
       LB2D_shift_0 <= LB2D_shift_0;
       LB2D_shift_1 <= LB2D_shift_1;
       LB2D_shift_2 <= LB2D_shift_2;
       LB2D_shift_3 <= LB2D_shift_3;
       LB2D_shift_4 <= LB2D_shift_4;
       LB2D_shift_5 <= LB2D_shift_5;
       LB2D_shift_6 <= LB2D_shift_6;
       LB2D_shift_7 <= LB2D_shift_7;
       LB2D_w_idx <= LB2D_w_idx;
       LB2D_x_idx <= LB2D_x_idx;
       LB2D_y_idx <= LB2D_y_idx;
       arg_0_TDATA <= arg_0_TDATA;
       arg_0_TVALID <= arg_0_TVALID;
       arg_1_TREADY <= arg_1_TREADY;
       slice_buff <= slice_buff;
       slice_full <= slice_full;
       stencil_buff <= stencil_buff;
       stencil_full <= stencil_full;
   end
   else if(step) begin
       LB2D_shift_0 <= n13;
       LB2D_shift_1 <= n16;
       LB2D_shift_2 <= n19;
       LB2D_shift_3 <= n22;
       LB2D_shift_4 <= n25;
       LB2D_shift_5 <= n28;
       LB2D_shift_6 <= n31;
       LB2D_shift_7 <= n34;
       LB2D_w_idx <= n42;
       LB2D_x_idx <= n48;
       LB2D_y_idx <= n55;
       arg_0_TDATA <= n58;
       arg_0_TVALID <= n61;
       arg_1_TREADY <= n64;
       slice_buff <= n148;
       slice_full <= n151;
       stencil_buff <= n315;
       stencil_full <= n318;
       LB2D_buff_0 [ LB2D_buff_0_addr0 ] <= LB2D_buff_0_data0;
       LB2D_buff_1 [ LB2D_buff_1_addr0 ] <= LB2D_buff_1_data0;
       LB2D_buff_2 [ LB2D_buff_2_addr0 ] <= LB2D_buff_2_data0;
       LB2D_buff_3 [ LB2D_buff_3_addr0 ] <= LB2D_buff_3_data0;
       LB2D_buff_4 [ LB2D_buff_4_addr0 ] <= LB2D_buff_4_data0;
       LB2D_buff_5 [ LB2D_buff_5_addr0 ] <= LB2D_buff_5_data0;
       LB2D_buff_6 [ LB2D_buff_6_addr0 ] <= LB2D_buff_6_data0;
       LB2D_buff_7 [ LB2D_buff_7_addr0 ] <= LB2D_buff_7_data0;
   end
end
endmodule
