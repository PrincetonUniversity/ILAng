module GB(
arg_0_TREADY,
arg_1_TDATA,
arg_1_TVALID,
RAM_w,
RAM_x,
RAM_y,
arg_0_TDATA,
arg_0_TVALID,
arg_1_TREADY,
cur_pix,
pre_pix,
proc_in,
st_ready,
stencil_0,
stencil_1,
stencil_2,
stencil_3,
stencil_4,
stencil_5,
stencil_6,
stencil_7,
stencil_8,
clk,rst,
step
);
input            arg_0_TREADY;
input      [7:0] arg_1_TDATA;
input            arg_1_TVALID;
input clk;
input rst;
input step;
output      [2:0] RAM_w;
output      [8:0] RAM_x;
output      [9:0] RAM_y;
output      [7:0] arg_0_TDATA;
output            arg_0_TVALID;
output            arg_1_TREADY;
output      [7:0] cur_pix;
output      [7:0] pre_pix;
output    [647:0] proc_in;
output            st_ready;
output     [71:0] stencil_0;
output     [71:0] stencil_1;
output     [71:0] stencil_2;
output     [71:0] stencil_3;
output     [71:0] stencil_4;
output     [71:0] stencil_5;
output     [71:0] stencil_6;
output     [71:0] stencil_7;
output     [71:0] stencil_8;
reg      [2:0] RAM_w;
reg      [8:0] RAM_x;
reg      [9:0] RAM_y;
reg      [7:0] arg_0_TDATA;
reg            arg_0_TVALID;
reg            arg_1_TREADY;
reg      [7:0] cur_pix;
reg      [7:0] pre_pix;
reg    [647:0] proc_in;
reg            st_ready;
reg     [71:0] stencil_0;
reg     [71:0] stencil_1;
reg     [71:0] stencil_2;
reg     [71:0] stencil_3;
reg     [71:0] stencil_4;
reg     [71:0] stencil_5;
reg     [71:0] stencil_6;
reg     [71:0] stencil_7;
reg     [71:0] stencil_8;
wire            arg_0_TREADY;
wire      [7:0] arg_1_TDATA;
wire            arg_1_TVALID;
wire            n0;
wire            n1;
wire            n2;
wire            n3;
wire            n4;
wire            n5;
wire            n6;
wire            n7;
wire            n8;
wire            n9;
wire            n10;
wire            n11;
wire            n12;
wire            n13;
wire      [2:0] n14;
wire      [2:0] n15;
wire      [2:0] n16;
wire            n17;
wire            n18;
wire            n19;
wire            n20;
wire      [2:0] n21;
wire      [2:0] n22;
wire      [2:0] n23;
wire      [8:0] n24;
wire      [8:0] n25;
wire      [8:0] n26;
wire      [8:0] n27;
wire      [8:0] n28;
wire            n29;
wire      [9:0] n30;
wire      [9:0] n31;
wire      [9:0] n32;
wire      [9:0] n33;
wire      [9:0] n34;
wire      [9:0] n35;
wire            n36;
wire      [7:0] n37;
wire      [7:0] n38;
wire      [7:0] n39;
wire      [7:0] n40;
wire      [7:0] n41;
wire      [7:0] n42;
wire      [7:0] n43;
wire      [7:0] n44;
wire      [7:0] n45;
wire     [15:0] n46;
wire     [23:0] n47;
wire     [31:0] n48;
wire     [39:0] n49;
wire     [47:0] n50;
wire     [55:0] n51;
wire     [63:0] n52;
wire     [71:0] n53;
wire      [7:0] n54;
wire      [7:0] n55;
wire      [7:0] n56;
wire      [7:0] n57;
wire      [7:0] n58;
wire      [7:0] n59;
wire      [7:0] n60;
wire      [7:0] n61;
wire      [7:0] n62;
wire     [15:0] n63;
wire     [23:0] n64;
wire     [31:0] n65;
wire     [39:0] n66;
wire     [47:0] n67;
wire     [55:0] n68;
wire     [63:0] n69;
wire     [71:0] n70;
wire      [7:0] n71;
wire      [7:0] n72;
wire      [7:0] n73;
wire      [7:0] n74;
wire      [7:0] n75;
wire      [7:0] n76;
wire      [7:0] n77;
wire      [7:0] n78;
wire      [7:0] n79;
wire     [15:0] n80;
wire     [23:0] n81;
wire     [31:0] n82;
wire     [39:0] n83;
wire     [47:0] n84;
wire     [55:0] n85;
wire     [63:0] n86;
wire     [71:0] n87;
wire      [7:0] n88;
wire      [7:0] n89;
wire      [7:0] n90;
wire      [7:0] n91;
wire      [7:0] n92;
wire      [7:0] n93;
wire      [7:0] n94;
wire      [7:0] n95;
wire      [7:0] n96;
wire     [15:0] n97;
wire     [23:0] n98;
wire     [31:0] n99;
wire     [39:0] n100;
wire     [47:0] n101;
wire     [55:0] n102;
wire     [63:0] n103;
wire     [71:0] n104;
wire      [7:0] n105;
wire      [7:0] n106;
wire      [7:0] n107;
wire      [7:0] n108;
wire      [7:0] n109;
wire      [7:0] n110;
wire      [7:0] n111;
wire      [7:0] n112;
wire      [7:0] n113;
wire     [15:0] n114;
wire     [23:0] n115;
wire     [31:0] n116;
wire     [39:0] n117;
wire     [47:0] n118;
wire     [55:0] n119;
wire     [63:0] n120;
wire     [71:0] n121;
wire      [7:0] n122;
wire      [7:0] n123;
wire      [7:0] n124;
wire      [7:0] n125;
wire      [7:0] n126;
wire      [7:0] n127;
wire      [7:0] n128;
wire      [7:0] n129;
wire      [7:0] n130;
wire     [15:0] n131;
wire     [23:0] n132;
wire     [31:0] n133;
wire     [39:0] n134;
wire     [47:0] n135;
wire     [55:0] n136;
wire     [63:0] n137;
wire     [71:0] n138;
wire      [7:0] n139;
wire      [7:0] n140;
wire      [7:0] n141;
wire      [7:0] n142;
wire      [7:0] n143;
wire      [7:0] n144;
wire      [7:0] n145;
wire      [7:0] n146;
wire      [7:0] n147;
wire     [15:0] n148;
wire     [23:0] n149;
wire     [31:0] n150;
wire     [39:0] n151;
wire     [47:0] n152;
wire     [55:0] n153;
wire     [63:0] n154;
wire     [71:0] n155;
wire      [7:0] n156;
wire      [7:0] n157;
wire      [7:0] n158;
wire      [7:0] n159;
wire      [7:0] n160;
wire      [7:0] n161;
wire      [7:0] n162;
wire      [7:0] n163;
wire      [7:0] n164;
wire     [15:0] n165;
wire     [23:0] n166;
wire     [31:0] n167;
wire     [39:0] n168;
wire     [47:0] n169;
wire     [55:0] n170;
wire     [63:0] n171;
wire     [71:0] n172;
wire      [7:0] n173;
wire      [7:0] n174;
wire      [7:0] n175;
wire      [7:0] n176;
wire      [7:0] n177;
wire      [7:0] n178;
wire      [7:0] n179;
wire      [7:0] n180;
wire      [7:0] n181;
wire     [15:0] n182;
wire     [23:0] n183;
wire     [31:0] n184;
wire     [39:0] n185;
wire     [47:0] n186;
wire     [55:0] n187;
wire     [63:0] n188;
wire     [71:0] n189;
wire    [143:0] n190;
wire    [215:0] n191;
wire    [287:0] n192;
wire    [359:0] n193;
wire    [431:0] n194;
wire    [503:0] n195;
wire    [575:0] n196;
wire    [647:0] n197;
wire    [647:0] n198;
wire      [7:0] n199;
wire      [7:0] n200;
wire      [7:0] n201;
wire      [7:0] n202;
wire            n203;
wire            n204;
wire            n205;
wire            n206;
wire            n207;
wire            n208;
wire            n209;
wire            n210;
wire            n211;
wire            n212;
wire            n213;
wire            n214;
wire            n215;
wire            n216;
wire      [7:0] n217;
wire      [7:0] n218;
wire      [7:0] n219;
wire      [7:0] n220;
wire      [7:0] n221;
wire    [647:0] n222;
wire    [647:0] n223;
wire            n224;
wire     [71:0] n225;
wire     [71:0] n226;
wire     [71:0] n227;
wire     [71:0] n228;
wire     [71:0] n229;
wire     [71:0] n230;
wire     [71:0] n231;
wire     [71:0] n232;
wire     [71:0] n233;
wire     [71:0] n234;
wire     [71:0] n235;
wire     [71:0] n236;
wire     [71:0] n237;
wire     [71:0] n238;
wire     [71:0] n239;
wire     [71:0] n240;
wire     [71:0] n241;
wire     [71:0] n242;
wire     [71:0] n243;
wire     [71:0] n244;
wire     [71:0] n245;
wire     [71:0] n246;
wire     [71:0] n247;
wire     [71:0] n248;
wire     [71:0] n249;
wire     [71:0] n250;
wire     [71:0] n251;
wire     [71:0] n252;
wire     [71:0] n253;
wire     [71:0] n254;
wire     [71:0] n255;
wire     [71:0] n256;
wire            n257;
wire      [8:0] n258;
wire      [7:0] n259;
wire            n260;
wire            n261;
wire            n262;
wire            n263;
wire            n264;
wire            n265;
wire      [7:0] n266;
wire      [7:0] n267;
wire      [7:0] n268;
wire      [7:0] n269;
wire      [7:0] n270;
wire      [7:0] n271;
wire      [7:0] n272;
wire      [7:0] n273;
wire      [7:0] n274;
wire      [7:0] n275;
wire      [7:0] n276;
wire      [7:0] n277;
wire      [7:0] n278;
wire      [7:0] n279;
wire      [7:0] n280;
wire      [7:0] n281;
wire      [7:0] n282;
wire      [7:0] n283;
wire      [7:0] n284;
wire      [7:0] n285;
wire      [7:0] n286;
wire      [7:0] n287;
wire      [7:0] n288;
wire      [7:0] n289;
wire      [7:0] n290;
wire      [7:0] n291;
wire      [7:0] n292;
wire      [7:0] n293;
wire      [7:0] n294;
wire      [7:0] n295;
wire      [7:0] n296;
wire      [7:0] n297;
wire      [7:0] n298;
wire      [7:0] n299;
wire      [7:0] n300;
wire      [7:0] n301;
wire      [7:0] n302;
wire      [7:0] n303;
wire      [7:0] n304;
wire      [7:0] n305;
wire      [7:0] n306;
wire      [7:0] n307;
wire      [7:0] n308;
wire      [7:0] n309;
wire      [7:0] n310;
wire      [7:0] n311;
wire      [7:0] n312;
wire      [7:0] n313;
wire      [7:0] n314;
wire      [7:0] n315;
wire      [7:0] n316;
wire      [7:0] n317;
wire      [7:0] n318;
wire      [7:0] n319;
wire      [7:0] n320;
wire      [7:0] n321;
wire      [7:0] n322;
wire      [7:0] n323;
wire      [7:0] n324;
wire      [7:0] n325;
wire      [7:0] n326;
wire      [7:0] n327;
wire      [7:0] n328;
wire     [15:0] n329;
wire     [23:0] n330;
wire     [31:0] n331;
wire     [39:0] n332;
wire     [47:0] n333;
wire     [55:0] n334;
wire     [63:0] n335;
wire     [71:0] n336;
wire     [71:0] n337;
wire     [71:0] n338;
wire     [71:0] n339;
wire     [71:0] n340;
wire      [8:0] RAM_0_addr0;
wire      [7:0] RAM_0_data0;
wire            n341;
wire            n342;
wire            n343;
wire            n344;
wire            n345;
wire            n346;
wire            n347;
wire            n348;
wire            n349;
wire            n350;
wire      [8:0] RAM_1_addr0;
wire      [7:0] RAM_1_data0;
wire            n351;
wire            n352;
wire            n353;
wire      [8:0] RAM_2_addr0;
wire      [7:0] RAM_2_data0;
wire            n354;
wire            n355;
wire            n356;
wire      [8:0] RAM_3_addr0;
wire      [7:0] RAM_3_data0;
wire            n357;
wire            n358;
wire            n359;
wire      [8:0] RAM_4_addr0;
wire      [7:0] RAM_4_data0;
wire            n360;
wire            n361;
wire            n362;
wire      [8:0] RAM_5_addr0;
wire      [7:0] RAM_5_data0;
wire            n363;
wire            n364;
wire            n365;
wire      [8:0] RAM_6_addr0;
wire      [7:0] RAM_6_data0;
wire            n366;
wire            n367;
wire            n368;
wire      [8:0] RAM_7_addr0;
wire      [7:0] RAM_7_data0;
wire            n369;
wire            n370;
wire            n371;
reg      [7:0] RAM_0[487:0];
reg      [7:0] RAM_1[487:0];
reg      [7:0] RAM_2[487:0];
reg      [7:0] RAM_3[487:0];
reg      [7:0] RAM_4[487:0];
reg      [7:0] RAM_5[487:0];
reg      [7:0] RAM_6[487:0];
reg      [7:0] RAM_7[487:0];
wire clk;
wire rst;
wire step;
assign n0 =  ( arg_1_TREADY ) == ( 1'd1 )  ;
assign n1 =  ( arg_0_TVALID ) == ( 1'd0 )  ;
assign n2 =  ( n0 ) & ( n1 )  ;
assign n3 =  ( arg_0_TREADY ) == ( 1'd0 )  ;
assign n4 =  ( n2 ) & ( n3 )  ;
assign n5 =  ( st_ready ) == ( 1'd0 )  ;
assign n6 =  ( n4 ) & ( n5 )  ;
assign n7 =  ( arg_1_TREADY ) == ( 1'd0 )  ;
assign n8 =  ( n7 ) & ( n1 )  ;
assign n9 =  ( n8 ) & ( n3 )  ;
assign n10 =  ( st_ready ) == ( 1'd1 )  ;
assign n11 =  ( n9 ) & ( n10 )  ;
assign n12 =  ( RAM_x ) == ( 9'd488 )  ;
assign n13 =  ( RAM_w ) == ( 3'd7 )  ;
assign n14 =  ( RAM_w ) + ( 3'd1 )  ;
assign n15 =  ( n13 ) ? ( 3'd0 ) : ( n14 ) ;
assign n16 =  ( n12 ) ? ( n15 ) : ( RAM_w ) ;
assign n17 =  ( arg_1_TVALID ) == ( 1'd1 )  ;
assign n18 =  ( n17 ) & ( n0 )  ;
assign n19 =  ( n18 ) & ( n1 )  ;
assign n20 =  ( n19 ) & ( n3 )  ;
assign n21 =  ( n20 ) ? ( RAM_w ) : ( RAM_w ) ;
assign n22 =  ( n11 ) ? ( n16 ) : ( n21 ) ;
assign n23 =  ( n6 ) ? ( RAM_w ) : ( n22 ) ;
assign n24 =  ( RAM_x ) + ( 9'd1 )  ;
assign n25 =  ( n12 ) ? ( 9'd1 ) : ( n24 ) ;
assign n26 =  ( n20 ) ? ( RAM_x ) : ( RAM_x ) ;
assign n27 =  ( n11 ) ? ( n25 ) : ( n26 ) ;
assign n28 =  ( n6 ) ? ( RAM_x ) : ( n27 ) ;
assign n29 =  ( RAM_y ) == ( 10'd648 )  ;
assign n30 =  ( RAM_y ) + ( 10'd1 )  ;
assign n31 =  ( n29 ) ? ( 10'd0 ) : ( n30 ) ;
assign n32 =  ( n12 ) ? ( n31 ) : ( RAM_y ) ;
assign n33 =  ( n20 ) ? ( RAM_y ) : ( RAM_y ) ;
assign n34 =  ( n11 ) ? ( n32 ) : ( n33 ) ;
assign n35 =  ( n6 ) ? ( RAM_y ) : ( n34 ) ;
assign n36 =  ( RAM_x ) > ( 9'd9 )  ;
assign n37 = stencil_8[71:64] ;
assign n38 = stencil_7[71:64] ;
assign n39 = stencil_6[71:64] ;
assign n40 = stencil_5[71:64] ;
assign n41 = stencil_4[71:64] ;
assign n42 = stencil_3[71:64] ;
assign n43 = stencil_2[71:64] ;
assign n44 = stencil_1[71:64] ;
assign n45 = stencil_0[71:64] ;
assign n46 =  { ( n44 ) , ( n45 ) }  ;
assign n47 =  { ( n43 ) , ( n46 ) }  ;
assign n48 =  { ( n42 ) , ( n47 ) }  ;
assign n49 =  { ( n41 ) , ( n48 ) }  ;
assign n50 =  { ( n40 ) , ( n49 ) }  ;
assign n51 =  { ( n39 ) , ( n50 ) }  ;
assign n52 =  { ( n38 ) , ( n51 ) }  ;
assign n53 =  { ( n37 ) , ( n52 ) }  ;
assign n54 = stencil_8[63:56] ;
assign n55 = stencil_7[63:56] ;
assign n56 = stencil_6[63:56] ;
assign n57 = stencil_5[63:56] ;
assign n58 = stencil_4[63:56] ;
assign n59 = stencil_3[63:56] ;
assign n60 = stencil_2[63:56] ;
assign n61 = stencil_1[63:56] ;
assign n62 = stencil_0[63:56] ;
assign n63 =  { ( n61 ) , ( n62 ) }  ;
assign n64 =  { ( n60 ) , ( n63 ) }  ;
assign n65 =  { ( n59 ) , ( n64 ) }  ;
assign n66 =  { ( n58 ) , ( n65 ) }  ;
assign n67 =  { ( n57 ) , ( n66 ) }  ;
assign n68 =  { ( n56 ) , ( n67 ) }  ;
assign n69 =  { ( n55 ) , ( n68 ) }  ;
assign n70 =  { ( n54 ) , ( n69 ) }  ;
assign n71 = stencil_8[55:48] ;
assign n72 = stencil_7[55:48] ;
assign n73 = stencil_6[55:48] ;
assign n74 = stencil_5[55:48] ;
assign n75 = stencil_4[55:48] ;
assign n76 = stencil_3[55:48] ;
assign n77 = stencil_2[55:48] ;
assign n78 = stencil_1[55:48] ;
assign n79 = stencil_0[55:48] ;
assign n80 =  { ( n78 ) , ( n79 ) }  ;
assign n81 =  { ( n77 ) , ( n80 ) }  ;
assign n82 =  { ( n76 ) , ( n81 ) }  ;
assign n83 =  { ( n75 ) , ( n82 ) }  ;
assign n84 =  { ( n74 ) , ( n83 ) }  ;
assign n85 =  { ( n73 ) , ( n84 ) }  ;
assign n86 =  { ( n72 ) , ( n85 ) }  ;
assign n87 =  { ( n71 ) , ( n86 ) }  ;
assign n88 = stencil_8[47:40] ;
assign n89 = stencil_7[47:40] ;
assign n90 = stencil_6[47:40] ;
assign n91 = stencil_5[47:40] ;
assign n92 = stencil_4[47:40] ;
assign n93 = stencil_3[47:40] ;
assign n94 = stencil_2[47:40] ;
assign n95 = stencil_1[47:40] ;
assign n96 = stencil_0[47:40] ;
assign n97 =  { ( n95 ) , ( n96 ) }  ;
assign n98 =  { ( n94 ) , ( n97 ) }  ;
assign n99 =  { ( n93 ) , ( n98 ) }  ;
assign n100 =  { ( n92 ) , ( n99 ) }  ;
assign n101 =  { ( n91 ) , ( n100 ) }  ;
assign n102 =  { ( n90 ) , ( n101 ) }  ;
assign n103 =  { ( n89 ) , ( n102 ) }  ;
assign n104 =  { ( n88 ) , ( n103 ) }  ;
assign n105 = stencil_8[39:32] ;
assign n106 = stencil_7[39:32] ;
assign n107 = stencil_6[39:32] ;
assign n108 = stencil_5[39:32] ;
assign n109 = stencil_4[39:32] ;
assign n110 = stencil_3[39:32] ;
assign n111 = stencil_2[39:32] ;
assign n112 = stencil_1[39:32] ;
assign n113 = stencil_0[39:32] ;
assign n114 =  { ( n112 ) , ( n113 ) }  ;
assign n115 =  { ( n111 ) , ( n114 ) }  ;
assign n116 =  { ( n110 ) , ( n115 ) }  ;
assign n117 =  { ( n109 ) , ( n116 ) }  ;
assign n118 =  { ( n108 ) , ( n117 ) }  ;
assign n119 =  { ( n107 ) , ( n118 ) }  ;
assign n120 =  { ( n106 ) , ( n119 ) }  ;
assign n121 =  { ( n105 ) , ( n120 ) }  ;
assign n122 = stencil_8[31:24] ;
assign n123 = stencil_7[31:24] ;
assign n124 = stencil_6[31:24] ;
assign n125 = stencil_5[31:24] ;
assign n126 = stencil_4[31:24] ;
assign n127 = stencil_3[31:24] ;
assign n128 = stencil_2[31:24] ;
assign n129 = stencil_1[31:24] ;
assign n130 = stencil_0[31:24] ;
assign n131 =  { ( n129 ) , ( n130 ) }  ;
assign n132 =  { ( n128 ) , ( n131 ) }  ;
assign n133 =  { ( n127 ) , ( n132 ) }  ;
assign n134 =  { ( n126 ) , ( n133 ) }  ;
assign n135 =  { ( n125 ) , ( n134 ) }  ;
assign n136 =  { ( n124 ) , ( n135 ) }  ;
assign n137 =  { ( n123 ) , ( n136 ) }  ;
assign n138 =  { ( n122 ) , ( n137 ) }  ;
assign n139 = stencil_8[23:16] ;
assign n140 = stencil_7[23:16] ;
assign n141 = stencil_6[23:16] ;
assign n142 = stencil_5[23:16] ;
assign n143 = stencil_4[23:16] ;
assign n144 = stencil_3[23:16] ;
assign n145 = stencil_2[23:16] ;
assign n146 = stencil_1[23:16] ;
assign n147 = stencil_0[23:16] ;
assign n148 =  { ( n146 ) , ( n147 ) }  ;
assign n149 =  { ( n145 ) , ( n148 ) }  ;
assign n150 =  { ( n144 ) , ( n149 ) }  ;
assign n151 =  { ( n143 ) , ( n150 ) }  ;
assign n152 =  { ( n142 ) , ( n151 ) }  ;
assign n153 =  { ( n141 ) , ( n152 ) }  ;
assign n154 =  { ( n140 ) , ( n153 ) }  ;
assign n155 =  { ( n139 ) , ( n154 ) }  ;
assign n156 = stencil_8[15:8] ;
assign n157 = stencil_7[15:8] ;
assign n158 = stencil_6[15:8] ;
assign n159 = stencil_5[15:8] ;
assign n160 = stencil_4[15:8] ;
assign n161 = stencil_3[15:8] ;
assign n162 = stencil_2[15:8] ;
assign n163 = stencil_1[15:8] ;
assign n164 = stencil_0[15:8] ;
assign n165 =  { ( n163 ) , ( n164 ) }  ;
assign n166 =  { ( n162 ) , ( n165 ) }  ;
assign n167 =  { ( n161 ) , ( n166 ) }  ;
assign n168 =  { ( n160 ) , ( n167 ) }  ;
assign n169 =  { ( n159 ) , ( n168 ) }  ;
assign n170 =  { ( n158 ) , ( n169 ) }  ;
assign n171 =  { ( n157 ) , ( n170 ) }  ;
assign n172 =  { ( n156 ) , ( n171 ) }  ;
assign n173 = stencil_8[7:0] ;
assign n174 = stencil_7[7:0] ;
assign n175 = stencil_6[7:0] ;
assign n176 = stencil_5[7:0] ;
assign n177 = stencil_4[7:0] ;
assign n178 = stencil_3[7:0] ;
assign n179 = stencil_2[7:0] ;
assign n180 = stencil_1[7:0] ;
assign n181 = stencil_0[7:0] ;
assign n182 =  { ( n180 ) , ( n181 ) }  ;
assign n183 =  { ( n179 ) , ( n182 ) }  ;
assign n184 =  { ( n178 ) , ( n183 ) }  ;
assign n185 =  { ( n177 ) , ( n184 ) }  ;
assign n186 =  { ( n176 ) , ( n185 ) }  ;
assign n187 =  { ( n175 ) , ( n186 ) }  ;
assign n188 =  { ( n174 ) , ( n187 ) }  ;
assign n189 =  { ( n173 ) , ( n188 ) }  ;
assign n190 =  { ( n172 ) , ( n189 ) }  ;
assign n191 =  { ( n155 ) , ( n190 ) }  ;
assign n192 =  { ( n138 ) , ( n191 ) }  ;
assign n193 =  { ( n121 ) , ( n192 ) }  ;
assign n194 =  { ( n104 ) , ( n193 ) }  ;
assign n195 =  { ( n87 ) , ( n194 ) }  ;
assign n196 =  { ( n70 ) , ( n195 ) }  ;
assign n197 =  { ( n53 ) , ( n196 ) }  ;
assign n198 =  ( n36 ) ? ( n197 ) : ( proc_in ) ;
//assign n199 = gb_fun(n198) ;
gb_fun gb_fun_U (
        .a (n198),
        .b (n199)
        );

assign n200 =  ( n20 ) ? ( arg_0_TDATA ) : ( arg_0_TDATA ) ;
assign n201 =  ( n11 ) ? ( arg_0_TDATA ) : ( n200 ) ;
assign n202 =  ( n6 ) ? ( n199 ) : ( n201 ) ;
assign n203 =  ( RAM_x ) > ( 9'd8 )  ;
assign n204 =  ( RAM_y ) >= ( 10'd8 )  ;
assign n205 =  ( n203 ) & ( n204 )  ;
assign n206 =  ( RAM_x ) == ( 9'd1 )  ;
assign n207 =  ( RAM_y ) > ( 10'd8 )  ;
assign n208 =  ( n206 ) & ( n207 )  ;
assign n209 =  ( n205 ) | ( n208 )  ;
assign n210 =  ( n209 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n211 =  ( n20 ) ? ( 1'd0 ) : ( arg_0_TVALID ) ;
assign n212 =  ( n11 ) ? ( 1'd0 ) : ( n211 ) ;
assign n213 =  ( n6 ) ? ( n210 ) : ( n212 ) ;
assign n214 =  ( n20 ) ? ( 1'd0 ) : ( arg_1_TREADY ) ;
assign n215 =  ( n11 ) ? ( 1'd1 ) : ( n214 ) ;
assign n216 =  ( n6 ) ? ( 1'd1 ) : ( n215 ) ;
assign n217 =  ( n20 ) ? ( arg_1_TDATA ) : ( cur_pix ) ;
assign n218 =  ( n11 ) ? ( n217 ) : ( n217 ) ;
assign n219 =  ( n6 ) ? ( cur_pix ) : ( n218 ) ;
assign n220 =  ( n11 ) ? ( cur_pix ) : ( pre_pix ) ;
assign n221 =  ( n6 ) ? ( pre_pix ) : ( n220 ) ;
assign n222 =  ( n11 ) ? ( proc_in ) : ( proc_in ) ;
assign n223 =  ( n6 ) ? ( n198 ) : ( n222 ) ;
assign n224 =  ( RAM_y ) < ( 10'd8 )  ;
assign n225 =  ( n224 ) ? ( stencil_0 ) : ( stencil_1 ) ;
assign n226 =  ( n20 ) ? ( stencil_0 ) : ( stencil_0 ) ;
assign n227 =  ( n11 ) ? ( stencil_0 ) : ( n226 ) ;
assign n228 =  ( n6 ) ? ( n225 ) : ( n227 ) ;
assign n229 =  ( n224 ) ? ( stencil_1 ) : ( stencil_2 ) ;
assign n230 =  ( n20 ) ? ( stencil_1 ) : ( stencil_1 ) ;
assign n231 =  ( n11 ) ? ( stencil_1 ) : ( n230 ) ;
assign n232 =  ( n6 ) ? ( n229 ) : ( n231 ) ;
assign n233 =  ( n224 ) ? ( stencil_2 ) : ( stencil_3 ) ;
assign n234 =  ( n20 ) ? ( stencil_2 ) : ( stencil_2 ) ;
assign n235 =  ( n11 ) ? ( stencil_2 ) : ( n234 ) ;
assign n236 =  ( n6 ) ? ( n233 ) : ( n235 ) ;
assign n237 =  ( n224 ) ? ( stencil_3 ) : ( stencil_4 ) ;
assign n238 =  ( n20 ) ? ( stencil_3 ) : ( stencil_3 ) ;
assign n239 =  ( n11 ) ? ( stencil_3 ) : ( n238 ) ;
assign n240 =  ( n6 ) ? ( n237 ) : ( n239 ) ;
assign n241 =  ( n224 ) ? ( stencil_4 ) : ( stencil_5 ) ;
assign n242 =  ( n20 ) ? ( stencil_4 ) : ( stencil_4 ) ;
assign n243 =  ( n11 ) ? ( stencil_4 ) : ( n242 ) ;
assign n244 =  ( n6 ) ? ( n241 ) : ( n243 ) ;
assign n245 =  ( n224 ) ? ( stencil_5 ) : ( stencil_6 ) ;
assign n246 =  ( n20 ) ? ( stencil_5 ) : ( stencil_5 ) ;
assign n247 =  ( n11 ) ? ( stencil_5 ) : ( n246 ) ;
assign n248 =  ( n6 ) ? ( n245 ) : ( n247 ) ;
assign n249 =  ( n224 ) ? ( stencil_6 ) : ( stencil_7 ) ;
assign n250 =  ( n20 ) ? ( stencil_6 ) : ( stencil_6 ) ;
assign n251 =  ( n11 ) ? ( stencil_6 ) : ( n250 ) ;
assign n252 =  ( n6 ) ? ( n249 ) : ( n251 ) ;
assign n253 =  ( n224 ) ? ( stencil_7 ) : ( stencil_8 ) ;
assign n254 =  ( n20 ) ? ( stencil_7 ) : ( stencil_7 ) ;
assign n255 =  ( n11 ) ? ( stencil_7 ) : ( n254 ) ;
assign n256 =  ( n6 ) ? ( n253 ) : ( n255 ) ;
assign n257 =  ( RAM_w ) == ( 3'd0 )  ;
assign n258 =  ( RAM_x ) - ( 9'd1 )  ;
assign n259 =  (  RAM_7 [ n258 ] )  ;
assign n260 =  ( RAM_w ) == ( 3'd1 )  ;
assign n261 =  ( RAM_w ) == ( 3'd2 )  ;
assign n262 =  ( RAM_w ) == ( 3'd3 )  ;
assign n263 =  ( RAM_w ) == ( 3'd4 )  ;
assign n264 =  ( RAM_w ) == ( 3'd5 )  ;
assign n265 =  ( RAM_w ) == ( 3'd6 )  ;
assign n266 =  (  RAM_6 [ n258 ] )  ;
assign n267 =  ( n265 ) ? ( n259 ) : ( n266 ) ;
assign n268 =  ( n264 ) ? ( n259 ) : ( n267 ) ;
assign n269 =  ( n263 ) ? ( n259 ) : ( n268 ) ;
assign n270 =  ( n262 ) ? ( n259 ) : ( n269 ) ;
assign n271 =  ( n261 ) ? ( n259 ) : ( n270 ) ;
assign n272 =  ( n260 ) ? ( n259 ) : ( n271 ) ;
assign n273 =  ( n257 ) ? ( n259 ) : ( n272 ) ;
assign n274 =  (  RAM_5 [ n258 ] )  ;
assign n275 =  ( n265 ) ? ( n266 ) : ( n274 ) ;
assign n276 =  ( n264 ) ? ( n266 ) : ( n275 ) ;
assign n277 =  ( n263 ) ? ( n266 ) : ( n276 ) ;
assign n278 =  ( n262 ) ? ( n266 ) : ( n277 ) ;
assign n279 =  ( n261 ) ? ( n266 ) : ( n278 ) ;
assign n280 =  ( n260 ) ? ( n266 ) : ( n279 ) ;
assign n281 =  ( n257 ) ? ( n266 ) : ( n280 ) ;
assign n282 =  (  RAM_4 [ n258 ] )  ;
assign n283 =  ( n265 ) ? ( n274 ) : ( n282 ) ;
assign n284 =  ( n264 ) ? ( n274 ) : ( n283 ) ;
assign n285 =  ( n263 ) ? ( n274 ) : ( n284 ) ;
assign n286 =  ( n262 ) ? ( n274 ) : ( n285 ) ;
assign n287 =  ( n261 ) ? ( n274 ) : ( n286 ) ;
assign n288 =  ( n260 ) ? ( n274 ) : ( n287 ) ;
assign n289 =  ( n257 ) ? ( n274 ) : ( n288 ) ;
assign n290 =  (  RAM_3 [ n258 ] )  ;
assign n291 =  ( n265 ) ? ( n282 ) : ( n290 ) ;
assign n292 =  ( n264 ) ? ( n282 ) : ( n291 ) ;
assign n293 =  ( n263 ) ? ( n282 ) : ( n292 ) ;
assign n294 =  ( n262 ) ? ( n282 ) : ( n293 ) ;
assign n295 =  ( n261 ) ? ( n282 ) : ( n294 ) ;
assign n296 =  ( n260 ) ? ( n282 ) : ( n295 ) ;
assign n297 =  ( n257 ) ? ( n282 ) : ( n296 ) ;
assign n298 =  (  RAM_2 [ n258 ] )  ;
assign n299 =  ( n265 ) ? ( n290 ) : ( n298 ) ;
assign n300 =  ( n264 ) ? ( n290 ) : ( n299 ) ;
assign n301 =  ( n263 ) ? ( n290 ) : ( n300 ) ;
assign n302 =  ( n262 ) ? ( n290 ) : ( n301 ) ;
assign n303 =  ( n261 ) ? ( n290 ) : ( n302 ) ;
assign n304 =  ( n260 ) ? ( n290 ) : ( n303 ) ;
assign n305 =  ( n257 ) ? ( n290 ) : ( n304 ) ;
assign n306 =  (  RAM_1 [ n258 ] )  ;
assign n307 =  ( n265 ) ? ( n298 ) : ( n306 ) ;
assign n308 =  ( n264 ) ? ( n298 ) : ( n307 ) ;
assign n309 =  ( n263 ) ? ( n298 ) : ( n308 ) ;
assign n310 =  ( n262 ) ? ( n298 ) : ( n309 ) ;
assign n311 =  ( n261 ) ? ( n298 ) : ( n310 ) ;
assign n312 =  ( n260 ) ? ( n298 ) : ( n311 ) ;
assign n313 =  ( n257 ) ? ( n298 ) : ( n312 ) ;
assign n314 =  (  RAM_0 [ n258 ] )  ;
assign n315 =  ( n265 ) ? ( n306 ) : ( n314 ) ;
assign n316 =  ( n264 ) ? ( n306 ) : ( n315 ) ;
assign n317 =  ( n263 ) ? ( n306 ) : ( n316 ) ;
assign n318 =  ( n262 ) ? ( n306 ) : ( n317 ) ;
assign n319 =  ( n261 ) ? ( n306 ) : ( n318 ) ;
assign n320 =  ( n260 ) ? ( n306 ) : ( n319 ) ;
assign n321 =  ( n257 ) ? ( n306 ) : ( n320 ) ;
assign n322 =  ( n265 ) ? ( n314 ) : ( n259 ) ;
assign n323 =  ( n264 ) ? ( n314 ) : ( n322 ) ;
assign n324 =  ( n263 ) ? ( n314 ) : ( n323 ) ;
assign n325 =  ( n262 ) ? ( n314 ) : ( n324 ) ;
assign n326 =  ( n261 ) ? ( n314 ) : ( n325 ) ;
assign n327 =  ( n260 ) ? ( n314 ) : ( n326 ) ;
assign n328 =  ( n257 ) ? ( n314 ) : ( n327 ) ;
assign n329 =  { ( n321 ) , ( n328 ) }  ;
assign n330 =  { ( n313 ) , ( n329 ) }  ;
assign n331 =  { ( n305 ) , ( n330 ) }  ;
assign n332 =  { ( n297 ) , ( n331 ) }  ;
assign n333 =  { ( n289 ) , ( n332 ) }  ;
assign n334 =  { ( n281 ) , ( n333 ) }  ;
assign n335 =  { ( n273 ) , ( n334 ) }  ;
assign n336 =  { ( pre_pix ) , ( n335 ) }  ;
assign n337 =  ( n224 ) ? ( stencil_8 ) : ( n336 ) ;
assign n338 =  ( n20 ) ? ( stencil_8 ) : ( stencil_8 ) ;
assign n339 =  ( n11 ) ? ( n337 ) : ( n338 ) ;
assign n340 =  ( n6 ) ? ( stencil_8 ) : ( n339 ) ;
assign n341 = ~ ( n6 ) ;
assign n342 = ~ ( n11 ) ;
assign n343 =  ( n341 ) & ( n342 )  ;
assign n344 = ~ ( n20 ) ;
assign n345 =  ( n343 ) & ( n344 )  ;
assign n346 =  ( n343 ) & ( n20 )  ;
assign n347 =  ( n341 ) & ( n11 )  ;
assign n348 = ~ ( n257 ) ;
assign n349 =  ( n347 ) & ( n348 )  ;
assign n350 =  ( n347 ) & ( n257 )  ;
assign RAM_0_addr0 = n350 ? (n258) : (0);
assign RAM_0_data0 = n350 ? (pre_pix) : (RAM_0[0]);
assign n351 = ~ ( n260 ) ;
assign n352 =  ( n347 ) & ( n351 )  ;
assign n353 =  ( n347 ) & ( n260 )  ;
assign RAM_1_addr0 = n353 ? (n258) : (0);
assign RAM_1_data0 = n353 ? (pre_pix) : (RAM_1[0]);
assign n354 = ~ ( n261 ) ;
assign n355 =  ( n347 ) & ( n354 )  ;
assign n356 =  ( n347 ) & ( n261 )  ;
assign RAM_2_addr0 = n356 ? (n258) : (0);
assign RAM_2_data0 = n356 ? (pre_pix) : (RAM_2[0]);
assign n357 = ~ ( n262 ) ;
assign n358 =  ( n347 ) & ( n357 )  ;
assign n359 =  ( n347 ) & ( n262 )  ;
assign RAM_3_addr0 = n359 ? (n258) : (0);
assign RAM_3_data0 = n359 ? (pre_pix) : (RAM_3[0]);
assign n360 = ~ ( n263 ) ;
assign n361 =  ( n347 ) & ( n360 )  ;
assign n362 =  ( n347 ) & ( n263 )  ;
assign RAM_4_addr0 = n362 ? (n258) : (0);
assign RAM_4_data0 = n362 ? (pre_pix) : (RAM_4[0]);
assign n363 = ~ ( n264 ) ;
assign n364 =  ( n347 ) & ( n363 )  ;
assign n365 =  ( n347 ) & ( n264 )  ;
assign RAM_5_addr0 = n365 ? (n258) : (0);
assign RAM_5_data0 = n365 ? (pre_pix) : (RAM_5[0]);
assign n366 = ~ ( n265 ) ;
assign n367 =  ( n347 ) & ( n366 )  ;
assign n368 =  ( n347 ) & ( n265 )  ;
assign RAM_6_addr0 = n368 ? (n258) : (0);
assign RAM_6_data0 = n368 ? (pre_pix) : (RAM_6[0]);
assign n369 = ~ ( n13 ) ;
assign n370 =  ( n347 ) & ( n369 )  ;
assign n371 =  ( n347 ) & ( n13 )  ;
assign RAM_7_addr0 = n371 ? (n258) : (0);
assign RAM_7_data0 = n371 ? (pre_pix) : (RAM_7[0]);
/*
function [7:0] gb_fun ;
input [647:0] arg0;
    begin
//TODO: Add the specific function HERE.    end
endfunction
*/

always @(posedge clk) begin
   if(rst) begin
       RAM_w <= RAM_w;
       RAM_x <= RAM_x;
       RAM_y <= RAM_y;
       arg_0_TDATA <= arg_0_TDATA;
       arg_0_TVALID <= arg_0_TVALID;
       arg_1_TREADY <= arg_1_TREADY;
       cur_pix <= cur_pix;
       pre_pix <= pre_pix;
       proc_in <= proc_in;
       st_ready <= st_ready;
       stencil_0 <= stencil_0;
       stencil_1 <= stencil_1;
       stencil_2 <= stencil_2;
       stencil_3 <= stencil_3;
       stencil_4 <= stencil_4;
       stencil_5 <= stencil_5;
       stencil_6 <= stencil_6;
       stencil_7 <= stencil_7;
       stencil_8 <= stencil_8;
   end
   else if(step) begin
       RAM_w <= n23;
       RAM_x <= n28;
       RAM_y <= n35;
       arg_0_TDATA <= n202;
       arg_0_TVALID <= n213;
       arg_1_TREADY <= n216;
       cur_pix <= n219;
       pre_pix <= n221;
       proc_in <= n223;
       st_ready <= st_ready;
       stencil_0 <= n228;
       stencil_1 <= n232;
       stencil_2 <= n236;
       stencil_3 <= n240;
       stencil_4 <= n244;
       stencil_5 <= n248;
       stencil_6 <= n252;
       stencil_7 <= n256;
       stencil_8 <= n340;
       RAM_0 [ RAM_0_addr0 ] <= RAM_0_data0;
       RAM_1 [ RAM_1_addr0 ] <= RAM_1_data0;
       RAM_2 [ RAM_2_addr0 ] <= RAM_2_data0;
       RAM_3 [ RAM_3_addr0 ] <= RAM_3_data0;
       RAM_4 [ RAM_4_addr0 ] <= RAM_4_data0;
       RAM_5 [ RAM_5_addr0 ] <= RAM_5_data0;
       RAM_6 [ RAM_6_addr0 ] <= RAM_6_data0;
       RAM_7 [ RAM_7_addr0 ] <= RAM_7_data0;
   end
end
endmodule
