module counter(input clk, input rst, input en, output reg full, inout p, inout q, output reg ro, output reg roi); // no semicolon

wire a;
reg b;
wire a;
reg b;

wire full;
wire p;

reg roi;

endmodule

