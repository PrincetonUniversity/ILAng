module SPEC_A(
arg_0_TREADY,
arg_1_TDATA,
arg_1_TVALID,
RAM_w,
RAM_x,
RAM_y,
arg_0_TDATA,
arg_0_TVALID,
arg_1_TREADY,
cur_pix,
gbit,
pre_pix,
proc_in,
st_ready,
stencil_0,
stencil_1,
stencil_2,
stencil_3,
stencil_4,
stencil_5,
stencil_6,
stencil_7,
stencil_8,
clk,rst,
step
);
input            arg_0_TREADY;
input      [7:0] arg_1_TDATA;
input            arg_1_TVALID;
input clk;
input rst;
input step;
output      [2:0] RAM_w;
output      [8:0] RAM_x;
output      [9:0] RAM_y;
output      [7:0] arg_0_TDATA;
output            arg_0_TVALID;
output            arg_1_TREADY;
output      [7:0] cur_pix;
output      [3:0] gbit;
output      [7:0] pre_pix;
output    [647:0] proc_in;
output            st_ready;
output     [71:0] stencil_0;
output     [71:0] stencil_1;
output     [71:0] stencil_2;
output     [71:0] stencil_3;
output     [71:0] stencil_4;
output     [71:0] stencil_5;
output     [71:0] stencil_6;
output     [71:0] stencil_7;
output     [71:0] stencil_8;
reg      [2:0] RAM_w;
reg      [8:0] RAM_x;
reg      [9:0] RAM_y;
reg      [7:0] arg_0_TDATA;
reg            arg_0_TVALID;
reg            arg_1_TREADY;
reg      [7:0] cur_pix;
reg      [3:0] gbit;
reg      [7:0] pre_pix;
reg    [647:0] proc_in;
reg            st_ready;
reg     [71:0] stencil_0;
reg     [71:0] stencil_1;
reg     [71:0] stencil_2;
reg     [71:0] stencil_3;
reg     [71:0] stencil_4;
reg     [71:0] stencil_5;
reg     [71:0] stencil_6;
reg     [71:0] stencil_7;
reg     [71:0] stencil_8;
wire            arg_0_TREADY;
wire      [7:0] arg_1_TDATA;
wire            arg_1_TVALID;
wire            n0;
wire            n1;
wire            n2;
wire            n3;
wire            n4;
wire            n5;
wire            n6;
wire            n7;
wire            n8;
wire            n9;
wire            n10;
wire            n11;
wire            n12;
wire            n13;
wire            n14;
wire            n15;
wire      [2:0] n16;
wire      [2:0] n17;
wire      [2:0] n18;
wire            n19;
wire            n20;
wire            n21;
wire            n22;
wire            n23;
wire            n24;
wire      [2:0] n25;
wire      [2:0] n26;
wire      [2:0] n27;
wire      [2:0] n28;
wire      [8:0] n29;
wire      [8:0] n30;
wire      [8:0] n31;
wire      [8:0] n32;
wire      [8:0] n33;
wire      [8:0] n34;
wire            n35;
wire      [9:0] n36;
wire      [9:0] n37;
wire      [9:0] n38;
wire      [9:0] n39;
wire      [9:0] n40;
wire      [9:0] n41;
wire      [9:0] n42;
wire            n43;
wire            n44;
wire            n45;
wire            n46;
wire            n47;
wire            n48;
wire            n49;
wire            n50;
wire      [7:0] n51;
wire      [7:0] n52;
wire      [7:0] n53;
wire      [7:0] n54;
wire      [7:0] n55;
wire      [7:0] n56;
wire      [7:0] n57;
wire      [7:0] n58;
wire      [7:0] n59;
wire     [15:0] n60;
wire     [23:0] n61;
wire     [31:0] n62;
wire     [39:0] n63;
wire     [47:0] n64;
wire     [55:0] n65;
wire     [63:0] n66;
wire     [71:0] n67;
wire      [7:0] n68;
wire      [7:0] n69;
wire      [7:0] n70;
wire      [7:0] n71;
wire      [7:0] n72;
wire      [7:0] n73;
wire      [7:0] n74;
wire      [7:0] n75;
wire      [7:0] n76;
wire     [15:0] n77;
wire     [23:0] n78;
wire     [31:0] n79;
wire     [39:0] n80;
wire     [47:0] n81;
wire     [55:0] n82;
wire     [63:0] n83;
wire     [71:0] n84;
wire      [7:0] n85;
wire      [7:0] n86;
wire      [7:0] n87;
wire      [7:0] n88;
wire      [7:0] n89;
wire      [7:0] n90;
wire      [7:0] n91;
wire      [7:0] n92;
wire      [7:0] n93;
wire     [15:0] n94;
wire     [23:0] n95;
wire     [31:0] n96;
wire     [39:0] n97;
wire     [47:0] n98;
wire     [55:0] n99;
wire     [63:0] n100;
wire     [71:0] n101;
wire      [7:0] n102;
wire      [7:0] n103;
wire      [7:0] n104;
wire      [7:0] n105;
wire      [7:0] n106;
wire      [7:0] n107;
wire      [7:0] n108;
wire      [7:0] n109;
wire      [7:0] n110;
wire     [15:0] n111;
wire     [23:0] n112;
wire     [31:0] n113;
wire     [39:0] n114;
wire     [47:0] n115;
wire     [55:0] n116;
wire     [63:0] n117;
wire     [71:0] n118;
wire      [7:0] n119;
wire      [7:0] n120;
wire      [7:0] n121;
wire      [7:0] n122;
wire      [7:0] n123;
wire      [7:0] n124;
wire      [7:0] n125;
wire      [7:0] n126;
wire      [7:0] n127;
wire     [15:0] n128;
wire     [23:0] n129;
wire     [31:0] n130;
wire     [39:0] n131;
wire     [47:0] n132;
wire     [55:0] n133;
wire     [63:0] n134;
wire     [71:0] n135;
wire      [7:0] n136;
wire      [7:0] n137;
wire      [7:0] n138;
wire      [7:0] n139;
wire      [7:0] n140;
wire      [7:0] n141;
wire      [7:0] n142;
wire      [7:0] n143;
wire      [7:0] n144;
wire     [15:0] n145;
wire     [23:0] n146;
wire     [31:0] n147;
wire     [39:0] n148;
wire     [47:0] n149;
wire     [55:0] n150;
wire     [63:0] n151;
wire     [71:0] n152;
wire      [7:0] n153;
wire      [7:0] n154;
wire      [7:0] n155;
wire      [7:0] n156;
wire      [7:0] n157;
wire      [7:0] n158;
wire      [7:0] n159;
wire      [7:0] n160;
wire      [7:0] n161;
wire     [15:0] n162;
wire     [23:0] n163;
wire     [31:0] n164;
wire     [39:0] n165;
wire     [47:0] n166;
wire     [55:0] n167;
wire     [63:0] n168;
wire     [71:0] n169;
wire      [7:0] n170;
wire      [7:0] n171;
wire      [7:0] n172;
wire      [7:0] n173;
wire      [7:0] n174;
wire      [7:0] n175;
wire      [7:0] n176;
wire      [7:0] n177;
wire      [7:0] n178;
wire     [15:0] n179;
wire     [23:0] n180;
wire     [31:0] n181;
wire     [39:0] n182;
wire     [47:0] n183;
wire     [55:0] n184;
wire     [63:0] n185;
wire     [71:0] n186;
wire      [7:0] n187;
wire      [7:0] n188;
wire      [7:0] n189;
wire      [7:0] n190;
wire      [7:0] n191;
wire      [7:0] n192;
wire      [7:0] n193;
wire      [7:0] n194;
wire      [7:0] n195;
wire     [15:0] n196;
wire     [23:0] n197;
wire     [31:0] n198;
wire     [39:0] n199;
wire     [47:0] n200;
wire     [55:0] n201;
wire     [63:0] n202;
wire     [71:0] n203;
wire    [143:0] n204;
wire    [215:0] n205;
wire    [287:0] n206;
wire    [359:0] n207;
wire    [431:0] n208;
wire    [503:0] n209;
wire    [575:0] n210;
wire    [647:0] n211;
wire    [647:0] n212;
wire    [647:0] n213;
wire      [7:0] n214;
wire      [7:0] n215;
wire      [7:0] n216;
wire      [7:0] n217;
wire      [7:0] n218;
wire      [7:0] n219;
wire            n220;
wire            n221;
wire            n222;
wire            n223;
wire            n224;
wire            n225;
wire      [8:0] n226;
wire            n227;
wire      [9:0] n228;
wire            n229;
wire            n230;
wire            n231;
wire            n232;
wire            n233;
wire            n234;
wire            n235;
wire            n236;
wire            n237;
wire      [7:0] n238;
wire      [7:0] n239;
wire      [7:0] n240;
wire      [7:0] n241;
wire      [7:0] n242;
wire      [7:0] n243;
wire      [7:0] n244;
wire    [647:0] n245;
wire    [647:0] n246;
wire    [647:0] n247;
wire            n248;
wire            n249;
wire            n250;
wire     [71:0] n251;
wire     [71:0] n252;
wire     [71:0] n253;
wire     [71:0] n254;
wire     [71:0] n255;
wire     [71:0] n256;
wire     [71:0] n257;
wire     [71:0] n258;
wire     [71:0] n259;
wire     [71:0] n260;
wire     [71:0] n261;
wire     [71:0] n262;
wire     [71:0] n263;
wire     [71:0] n264;
wire     [71:0] n265;
wire     [71:0] n266;
wire     [71:0] n267;
wire     [71:0] n268;
wire     [71:0] n269;
wire     [71:0] n270;
wire     [71:0] n271;
wire     [71:0] n272;
wire     [71:0] n273;
wire     [71:0] n274;
wire     [71:0] n275;
wire     [71:0] n276;
wire     [71:0] n277;
wire     [71:0] n278;
wire     [71:0] n279;
wire     [71:0] n280;
wire     [71:0] n281;
wire     [71:0] n282;
wire     [71:0] n283;
wire     [71:0] n284;
wire     [71:0] n285;
wire     [71:0] n286;
wire     [71:0] n287;
wire     [71:0] n288;
wire     [71:0] n289;
wire     [71:0] n290;
wire            n291;
wire      [8:0] n292;
wire      [7:0] n293;
wire            n294;
wire      [7:0] n295;
wire            n296;
wire      [7:0] n297;
wire            n298;
wire      [7:0] n299;
wire            n300;
wire      [7:0] n301;
wire            n302;
wire      [7:0] n303;
wire            n304;
wire      [7:0] n305;
wire      [7:0] n306;
wire      [7:0] n307;
wire      [7:0] n308;
wire      [7:0] n309;
wire      [7:0] n310;
wire      [7:0] n311;
wire      [7:0] n312;
wire      [7:0] n313;
wire      [7:0] n314;
wire      [7:0] n315;
wire      [7:0] n316;
wire      [7:0] n317;
wire      [7:0] n318;
wire      [7:0] n319;
wire      [7:0] n320;
wire      [7:0] n321;
wire      [7:0] n322;
wire      [7:0] n323;
wire      [7:0] n324;
wire      [7:0] n325;
wire      [7:0] n326;
wire      [7:0] n327;
wire      [7:0] n328;
wire      [7:0] n329;
wire      [7:0] n330;
wire      [7:0] n331;
wire      [7:0] n332;
wire      [7:0] n333;
wire      [7:0] n334;
wire      [7:0] n335;
wire      [7:0] n336;
wire      [7:0] n337;
wire      [7:0] n338;
wire      [7:0] n339;
wire      [7:0] n340;
wire      [7:0] n341;
wire      [7:0] n342;
wire      [7:0] n343;
wire      [7:0] n344;
wire      [7:0] n345;
wire      [7:0] n346;
wire      [7:0] n347;
wire      [7:0] n348;
wire      [7:0] n349;
wire      [7:0] n350;
wire      [7:0] n351;
wire      [7:0] n352;
wire      [7:0] n353;
wire      [7:0] n354;
wire      [7:0] n355;
wire      [7:0] n356;
wire      [7:0] n357;
wire      [7:0] n358;
wire      [7:0] n359;
wire      [7:0] n360;
wire      [7:0] n361;
wire      [7:0] n362;
wire     [15:0] n363;
wire     [23:0] n364;
wire     [31:0] n365;
wire     [39:0] n366;
wire     [47:0] n367;
wire     [55:0] n368;
wire     [63:0] n369;
wire     [71:0] n370;
wire     [71:0] n371;
wire     [71:0] n372;
wire     [71:0] n373;
wire     [71:0] n374;
wire     [71:0] n375;
wire      [8:0] RAM_0_addr0;
wire      [7:0] RAM_0_data0;
wire            n376;
wire            n377;
wire            n378;
wire            n379;
wire            n380;
wire            n381;
wire            n382;
wire            n383;
wire            n384;
wire            n385;
wire            n386;
wire            n387;
wire            n388;
wire      [8:0] RAM_1_addr0;
wire      [7:0] RAM_1_data0;
wire            n389;
wire            n390;
wire            n391;
wire      [8:0] RAM_2_addr0;
wire      [7:0] RAM_2_data0;
wire            n392;
wire            n393;
wire            n394;
wire      [8:0] RAM_3_addr0;
wire      [7:0] RAM_3_data0;
wire            n395;
wire            n396;
wire            n397;
wire      [8:0] RAM_4_addr0;
wire      [7:0] RAM_4_data0;
wire            n398;
wire            n399;
wire            n400;
wire      [8:0] RAM_5_addr0;
wire      [7:0] RAM_5_data0;
wire            n401;
wire            n402;
wire            n403;
wire      [8:0] RAM_6_addr0;
wire      [7:0] RAM_6_data0;
wire            n404;
wire            n405;
wire            n406;
wire      [8:0] RAM_7_addr0;
wire      [7:0] RAM_7_data0;
wire            n407;
wire            n408;
wire            n409;
reg      [7:0] RAM_0[487:0];
reg      [7:0] RAM_1[487:0];
reg      [7:0] RAM_2[487:0];
reg      [7:0] RAM_3[487:0];
reg      [7:0] RAM_4[487:0];
reg      [7:0] RAM_5[487:0];
reg      [7:0] RAM_6[487:0];
reg      [7:0] RAM_7[487:0];
wire clk;
wire rst;
wire step;
assign n0 =  ( arg_1_TREADY ) == ( 1'd0 )  ;
assign n1 =  ( arg_0_TREADY ) == ( 1'd0 )  ;
assign n2 =  ( n0 ) & ( n1 )  ;
assign n3 =  ( st_ready ) == ( 1'd0 )  ;
assign n4 =  ( n2 ) & ( n3 )  ;
assign n5 =  ( st_ready ) == ( 1'd1 )  ;
assign n6 =  ( n2 ) & ( n5 )  ;
assign n7 =  ( RAM_x ) == ( 9'd0 )  ;
assign n8 =  ( n6 ) & ( n7 )  ;
assign n9 =  ( RAM_y ) == ( 10'd0 )  ;
assign n10 =  ( n8 ) & ( n9 )  ;
assign n11 =  ( n7 ) & ( n9 )  ;
assign n12 = ~ ( n11 ) ;
assign n13 =  ( n6 ) & ( n12 )  ;
assign n14 =  ( RAM_x ) == ( 9'd488 )  ;
assign n15 =  ( RAM_w ) == ( 3'd7 )  ;
assign n16 =  ( RAM_w ) + ( 3'd1 )  ;
assign n17 =  ( n15 ) ? ( 3'd0 ) : ( n16 ) ;
assign n18 =  ( n14 ) ? ( n17 ) : ( RAM_w ) ;
assign n19 =  ( arg_1_TVALID ) == ( 1'd1 )  ;
assign n20 =  ( arg_1_TREADY ) == ( 1'd1 )  ;
assign n21 =  ( n19 ) & ( n20 )  ;
assign n22 =  ( arg_0_TVALID ) == ( 1'd0 )  ;
assign n23 =  ( n21 ) & ( n22 )  ;
assign n24 =  ( n23 ) & ( n1 )  ;
assign n25 =  ( n24 ) ? ( RAM_w ) : ( RAM_w ) ;
assign n26 =  ( n13 ) ? ( n18 ) : ( n25 ) ;
assign n27 =  ( n10 ) ? ( RAM_w ) : ( n26 ) ;
assign n28 =  ( n4 ) ? ( RAM_w ) : ( n27 ) ;
assign n29 =  ( RAM_x ) + ( 9'd1 )  ;
assign n30 =  ( n14 ) ? ( 9'd1 ) : ( n29 ) ;
assign n31 =  ( n24 ) ? ( RAM_x ) : ( RAM_x ) ;
assign n32 =  ( n13 ) ? ( n30 ) : ( n31 ) ;
assign n33 =  ( n10 ) ? ( 9'd1 ) : ( n32 ) ;
assign n34 =  ( n4 ) ? ( RAM_x ) : ( n33 ) ;
assign n35 =  ( RAM_y ) == ( 10'd648 )  ;
assign n36 =  ( RAM_y ) + ( 10'd1 )  ;
assign n37 =  ( n35 ) ? ( 10'd0 ) : ( n36 ) ;
assign n38 =  ( n14 ) ? ( n37 ) : ( RAM_y ) ;
assign n39 =  ( n24 ) ? ( RAM_y ) : ( RAM_y ) ;
assign n40 =  ( n13 ) ? ( n38 ) : ( n39 ) ;
assign n41 =  ( n10 ) ? ( RAM_y ) : ( n40 ) ;
assign n42 =  ( n4 ) ? ( RAM_y ) : ( n41 ) ;
assign n43 =  ( RAM_x ) == ( 9'd1 )  ;
assign n44 =  ( n43 ) & ( n35 )  ;
assign n45 =  ( RAM_x ) > ( 9'd8 )  ;
assign n46 =  ( RAM_y ) >= ( 10'd8 )  ;
assign n47 =  ( n45 ) & ( n46 )  ;
assign n48 =  ( RAM_y ) > ( 10'd8 )  ;
assign n49 =  ( n43 ) & ( n48 )  ;
assign n50 =  ( n47 ) | ( n49 )  ;
assign n51 = stencil_8[71:64] ;
assign n52 = stencil_7[71:64] ;
assign n53 = stencil_6[71:64] ;
assign n54 = stencil_5[71:64] ;
assign n55 = stencil_4[71:64] ;
assign n56 = stencil_3[71:64] ;
assign n57 = stencil_2[71:64] ;
assign n58 = stencil_1[71:64] ;
assign n59 = stencil_0[71:64] ;
assign n60 =  { ( n58 ) , ( n59 ) }  ;
assign n61 =  { ( n57 ) , ( n60 ) }  ;
assign n62 =  { ( n56 ) , ( n61 ) }  ;
assign n63 =  { ( n55 ) , ( n62 ) }  ;
assign n64 =  { ( n54 ) , ( n63 ) }  ;
assign n65 =  { ( n53 ) , ( n64 ) }  ;
assign n66 =  { ( n52 ) , ( n65 ) }  ;
assign n67 =  { ( n51 ) , ( n66 ) }  ;
assign n68 = stencil_8[63:56] ;
assign n69 = stencil_7[63:56] ;
assign n70 = stencil_6[63:56] ;
assign n71 = stencil_5[63:56] ;
assign n72 = stencil_4[63:56] ;
assign n73 = stencil_3[63:56] ;
assign n74 = stencil_2[63:56] ;
assign n75 = stencil_1[63:56] ;
assign n76 = stencil_0[63:56] ;
assign n77 =  { ( n75 ) , ( n76 ) }  ;
assign n78 =  { ( n74 ) , ( n77 ) }  ;
assign n79 =  { ( n73 ) , ( n78 ) }  ;
assign n80 =  { ( n72 ) , ( n79 ) }  ;
assign n81 =  { ( n71 ) , ( n80 ) }  ;
assign n82 =  { ( n70 ) , ( n81 ) }  ;
assign n83 =  { ( n69 ) , ( n82 ) }  ;
assign n84 =  { ( n68 ) , ( n83 ) }  ;
assign n85 = stencil_8[55:48] ;
assign n86 = stencil_7[55:48] ;
assign n87 = stencil_6[55:48] ;
assign n88 = stencil_5[55:48] ;
assign n89 = stencil_4[55:48] ;
assign n90 = stencil_3[55:48] ;
assign n91 = stencil_2[55:48] ;
assign n92 = stencil_1[55:48] ;
assign n93 = stencil_0[55:48] ;
assign n94 =  { ( n92 ) , ( n93 ) }  ;
assign n95 =  { ( n91 ) , ( n94 ) }  ;
assign n96 =  { ( n90 ) , ( n95 ) }  ;
assign n97 =  { ( n89 ) , ( n96 ) }  ;
assign n98 =  { ( n88 ) , ( n97 ) }  ;
assign n99 =  { ( n87 ) , ( n98 ) }  ;
assign n100 =  { ( n86 ) , ( n99 ) }  ;
assign n101 =  { ( n85 ) , ( n100 ) }  ;
assign n102 = stencil_8[47:40] ;
assign n103 = stencil_7[47:40] ;
assign n104 = stencil_6[47:40] ;
assign n105 = stencil_5[47:40] ;
assign n106 = stencil_4[47:40] ;
assign n107 = stencil_3[47:40] ;
assign n108 = stencil_2[47:40] ;
assign n109 = stencil_1[47:40] ;
assign n110 = stencil_0[47:40] ;
assign n111 =  { ( n109 ) , ( n110 ) }  ;
assign n112 =  { ( n108 ) , ( n111 ) }  ;
assign n113 =  { ( n107 ) , ( n112 ) }  ;
assign n114 =  { ( n106 ) , ( n113 ) }  ;
assign n115 =  { ( n105 ) , ( n114 ) }  ;
assign n116 =  { ( n104 ) , ( n115 ) }  ;
assign n117 =  { ( n103 ) , ( n116 ) }  ;
assign n118 =  { ( n102 ) , ( n117 ) }  ;
assign n119 = stencil_8[39:32] ;
assign n120 = stencil_7[39:32] ;
assign n121 = stencil_6[39:32] ;
assign n122 = stencil_5[39:32] ;
assign n123 = stencil_4[39:32] ;
assign n124 = stencil_3[39:32] ;
assign n125 = stencil_2[39:32] ;
assign n126 = stencil_1[39:32] ;
assign n127 = stencil_0[39:32] ;
assign n128 =  { ( n126 ) , ( n127 ) }  ;
assign n129 =  { ( n125 ) , ( n128 ) }  ;
assign n130 =  { ( n124 ) , ( n129 ) }  ;
assign n131 =  { ( n123 ) , ( n130 ) }  ;
assign n132 =  { ( n122 ) , ( n131 ) }  ;
assign n133 =  { ( n121 ) , ( n132 ) }  ;
assign n134 =  { ( n120 ) , ( n133 ) }  ;
assign n135 =  { ( n119 ) , ( n134 ) }  ;
assign n136 = stencil_8[31:24] ;
assign n137 = stencil_7[31:24] ;
assign n138 = stencil_6[31:24] ;
assign n139 = stencil_5[31:24] ;
assign n140 = stencil_4[31:24] ;
assign n141 = stencil_3[31:24] ;
assign n142 = stencil_2[31:24] ;
assign n143 = stencil_1[31:24] ;
assign n144 = stencil_0[31:24] ;
assign n145 =  { ( n143 ) , ( n144 ) }  ;
assign n146 =  { ( n142 ) , ( n145 ) }  ;
assign n147 =  { ( n141 ) , ( n146 ) }  ;
assign n148 =  { ( n140 ) , ( n147 ) }  ;
assign n149 =  { ( n139 ) , ( n148 ) }  ;
assign n150 =  { ( n138 ) , ( n149 ) }  ;
assign n151 =  { ( n137 ) , ( n150 ) }  ;
assign n152 =  { ( n136 ) , ( n151 ) }  ;
assign n153 = stencil_8[23:16] ;
assign n154 = stencil_7[23:16] ;
assign n155 = stencil_6[23:16] ;
assign n156 = stencil_5[23:16] ;
assign n157 = stencil_4[23:16] ;
assign n158 = stencil_3[23:16] ;
assign n159 = stencil_2[23:16] ;
assign n160 = stencil_1[23:16] ;
assign n161 = stencil_0[23:16] ;
assign n162 =  { ( n160 ) , ( n161 ) }  ;
assign n163 =  { ( n159 ) , ( n162 ) }  ;
assign n164 =  { ( n158 ) , ( n163 ) }  ;
assign n165 =  { ( n157 ) , ( n164 ) }  ;
assign n166 =  { ( n156 ) , ( n165 ) }  ;
assign n167 =  { ( n155 ) , ( n166 ) }  ;
assign n168 =  { ( n154 ) , ( n167 ) }  ;
assign n169 =  { ( n153 ) , ( n168 ) }  ;
assign n170 = stencil_8[15:8] ;
assign n171 = stencil_7[15:8] ;
assign n172 = stencil_6[15:8] ;
assign n173 = stencil_5[15:8] ;
assign n174 = stencil_4[15:8] ;
assign n175 = stencil_3[15:8] ;
assign n176 = stencil_2[15:8] ;
assign n177 = stencil_1[15:8] ;
assign n178 = stencil_0[15:8] ;
assign n179 =  { ( n177 ) , ( n178 ) }  ;
assign n180 =  { ( n176 ) , ( n179 ) }  ;
assign n181 =  { ( n175 ) , ( n180 ) }  ;
assign n182 =  { ( n174 ) , ( n181 ) }  ;
assign n183 =  { ( n173 ) , ( n182 ) }  ;
assign n184 =  { ( n172 ) , ( n183 ) }  ;
assign n185 =  { ( n171 ) , ( n184 ) }  ;
assign n186 =  { ( n170 ) , ( n185 ) }  ;
assign n187 = stencil_8[7:0] ;
assign n188 = stencil_7[7:0] ;
assign n189 = stencil_6[7:0] ;
assign n190 = stencil_5[7:0] ;
assign n191 = stencil_4[7:0] ;
assign n192 = stencil_3[7:0] ;
assign n193 = stencil_2[7:0] ;
assign n194 = stencil_1[7:0] ;
assign n195 = stencil_0[7:0] ;
assign n196 =  { ( n194 ) , ( n195 ) }  ;
assign n197 =  { ( n193 ) , ( n196 ) }  ;
assign n198 =  { ( n192 ) , ( n197 ) }  ;
assign n199 =  { ( n191 ) , ( n198 ) }  ;
assign n200 =  { ( n190 ) , ( n199 ) }  ;
assign n201 =  { ( n189 ) , ( n200 ) }  ;
assign n202 =  { ( n188 ) , ( n201 ) }  ;
assign n203 =  { ( n187 ) , ( n202 ) }  ;
assign n204 =  { ( n186 ) , ( n203 ) }  ;
assign n205 =  { ( n169 ) , ( n204 ) }  ;
assign n206 =  { ( n152 ) , ( n205 ) }  ;
assign n207 =  { ( n135 ) , ( n206 ) }  ;
assign n208 =  { ( n118 ) , ( n207 ) }  ;
assign n209 =  { ( n101 ) , ( n208 ) }  ;
assign n210 =  { ( n84 ) , ( n209 ) }  ;
assign n211 =  { ( n67 ) , ( n210 ) }  ;
assign n212 =  ( n50 ) ? ( n211 ) : ( proc_in ) ;
assign n213 =  ( n44 ) ? ( proc_in ) : ( n212 ) ;
//assign n214 = gb_fun(n213) ;
gb_fun gb_fun_U (
        .a (n213),
        .b (n214)
        );

assign n215 =  ( n44 ) ? ( arg_0_TDATA ) : ( n214 ) ;
assign n216 =  ( n24 ) ? ( arg_0_TDATA ) : ( arg_0_TDATA ) ;
assign n217 =  ( n13 ) ? ( arg_0_TDATA ) : ( n216 ) ;
assign n218 =  ( n10 ) ? ( arg_0_TDATA ) : ( n217 ) ;
assign n219 =  ( n4 ) ? ( n215 ) : ( n218 ) ;
assign n220 =  ( n50 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n221 =  ( n44 ) ? ( arg_0_TVALID ) : ( n220 ) ;
assign n222 =  ( n24 ) ? ( 1'd0 ) : ( arg_0_TVALID ) ;
assign n223 =  ( n13 ) ? ( arg_0_TVALID ) : ( n222 ) ;
assign n224 =  ( n10 ) ? ( 1'd0 ) : ( n223 ) ;
assign n225 =  ( n4 ) ? ( n221 ) : ( n224 ) ;
assign n226 =  ( 9'd488 ) - ( 9'd1 )  ;
assign n227 =  ( RAM_x ) == ( n226 )  ;
assign n228 =  ( 10'd648 ) - ( 10'd1 )  ;
assign n229 =  ( RAM_y ) == ( n228 )  ;
assign n230 =  ( n227 ) & ( n229 )  ;
assign n231 =  ( n230 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n232 =  ( RAM_y ) < ( 10'd8 )  ;
assign n233 =  ( n232 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n234 =  ( n24 ) ? ( 1'd0 ) : ( arg_1_TREADY ) ;
assign n235 =  ( n13 ) ? ( n233 ) : ( n234 ) ;
assign n236 =  ( n10 ) ? ( 1'd1 ) : ( n235 ) ;
assign n237 =  ( n4 ) ? ( n231 ) : ( n236 ) ;
assign n238 =  ( n24 ) ? ( arg_1_TDATA ) : ( cur_pix ) ;
assign n239 =  ( n13 ) ? ( cur_pix ) : ( n238 ) ;
assign n240 =  ( n10 ) ? ( cur_pix ) : ( n239 ) ;
assign n241 =  ( n4 ) ? ( cur_pix ) : ( n240 ) ;
assign n242 =  ( n13 ) ? ( cur_pix ) : ( pre_pix ) ;
assign n243 =  ( n10 ) ? ( cur_pix ) : ( n242 ) ;
assign n244 =  ( n4 ) ? ( pre_pix ) : ( n243 ) ;
assign n245 =  ( n13 ) ? ( proc_in ) : ( proc_in ) ;
assign n246 =  ( n10 ) ? ( proc_in ) : ( n245 ) ;
assign n247 =  ( n4 ) ? ( n213 ) : ( n246 ) ;
assign n248 =  ( n13 ) ? ( n233 ) : ( st_ready ) ;
assign n249 =  ( n10 ) ? ( 1'd1 ) : ( n248 ) ;
assign n250 =  ( n4 ) ? ( 1'd1 ) : ( n249 ) ;
assign n251 =  ( n232 ) ? ( stencil_0 ) : ( stencil_1 ) ;
assign n252 =  ( n24 ) ? ( stencil_0 ) : ( stencil_0 ) ;
assign n253 =  ( n13 ) ? ( stencil_0 ) : ( n252 ) ;
assign n254 =  ( n10 ) ? ( stencil_0 ) : ( n253 ) ;
assign n255 =  ( n4 ) ? ( n251 ) : ( n254 ) ;
assign n256 =  ( n232 ) ? ( stencil_1 ) : ( stencil_2 ) ;
assign n257 =  ( n24 ) ? ( stencil_1 ) : ( stencil_1 ) ;
assign n258 =  ( n13 ) ? ( stencil_1 ) : ( n257 ) ;
assign n259 =  ( n10 ) ? ( stencil_1 ) : ( n258 ) ;
assign n260 =  ( n4 ) ? ( n256 ) : ( n259 ) ;
assign n261 =  ( n232 ) ? ( stencil_2 ) : ( stencil_3 ) ;
assign n262 =  ( n24 ) ? ( stencil_2 ) : ( stencil_2 ) ;
assign n263 =  ( n13 ) ? ( stencil_2 ) : ( n262 ) ;
assign n264 =  ( n10 ) ? ( stencil_2 ) : ( n263 ) ;
assign n265 =  ( n4 ) ? ( n261 ) : ( n264 ) ;
assign n266 =  ( n232 ) ? ( stencil_3 ) : ( stencil_4 ) ;
assign n267 =  ( n24 ) ? ( stencil_3 ) : ( stencil_3 ) ;
assign n268 =  ( n13 ) ? ( stencil_3 ) : ( n267 ) ;
assign n269 =  ( n10 ) ? ( stencil_3 ) : ( n268 ) ;
assign n270 =  ( n4 ) ? ( n266 ) : ( n269 ) ;
assign n271 =  ( n232 ) ? ( stencil_4 ) : ( stencil_5 ) ;
assign n272 =  ( n24 ) ? ( stencil_4 ) : ( stencil_4 ) ;
assign n273 =  ( n13 ) ? ( stencil_4 ) : ( n272 ) ;
assign n274 =  ( n10 ) ? ( stencil_4 ) : ( n273 ) ;
assign n275 =  ( n4 ) ? ( n271 ) : ( n274 ) ;
assign n276 =  ( n232 ) ? ( stencil_5 ) : ( stencil_6 ) ;
assign n277 =  ( n24 ) ? ( stencil_5 ) : ( stencil_5 ) ;
assign n278 =  ( n13 ) ? ( stencil_5 ) : ( n277 ) ;
assign n279 =  ( n10 ) ? ( stencil_5 ) : ( n278 ) ;
assign n280 =  ( n4 ) ? ( n276 ) : ( n279 ) ;
assign n281 =  ( n232 ) ? ( stencil_6 ) : ( stencil_7 ) ;
assign n282 =  ( n24 ) ? ( stencil_6 ) : ( stencil_6 ) ;
assign n283 =  ( n13 ) ? ( stencil_6 ) : ( n282 ) ;
assign n284 =  ( n10 ) ? ( stencil_6 ) : ( n283 ) ;
assign n285 =  ( n4 ) ? ( n281 ) : ( n284 ) ;
assign n286 =  ( n232 ) ? ( stencil_7 ) : ( stencil_8 ) ;
assign n287 =  ( n24 ) ? ( stencil_7 ) : ( stencil_7 ) ;
assign n288 =  ( n13 ) ? ( stencil_7 ) : ( n287 ) ;
assign n289 =  ( n10 ) ? ( stencil_7 ) : ( n288 ) ;
assign n290 =  ( n4 ) ? ( n286 ) : ( n289 ) ;
assign n291 =  ( RAM_w ) == ( 3'd0 )  ;
assign n292 =  ( RAM_x ) - ( 9'd1 )  ;
assign n293 =  (  RAM_7 [ n292 ] )  ;
assign n294 =  ( RAM_w ) == ( 3'd1 )  ;
assign n295 =  (  RAM_0 [ n292 ] )  ;
assign n296 =  ( RAM_w ) == ( 3'd2 )  ;
assign n297 =  (  RAM_1 [ n292 ] )  ;
assign n298 =  ( RAM_w ) == ( 3'd3 )  ;
assign n299 =  (  RAM_2 [ n292 ] )  ;
assign n300 =  ( RAM_w ) == ( 3'd4 )  ;
assign n301 =  (  RAM_3 [ n292 ] )  ;
assign n302 =  ( RAM_w ) == ( 3'd5 )  ;
assign n303 =  (  RAM_4 [ n292 ] )  ;
assign n304 =  ( RAM_w ) == ( 3'd6 )  ;
assign n305 =  (  RAM_5 [ n292 ] )  ;
assign n306 =  (  RAM_6 [ n292 ] )  ;
assign n307 =  ( n304 ) ? ( n305 ) : ( n306 ) ;
assign n308 =  ( n302 ) ? ( n303 ) : ( n307 ) ;
assign n309 =  ( n300 ) ? ( n301 ) : ( n308 ) ;
assign n310 =  ( n298 ) ? ( n299 ) : ( n309 ) ;
assign n311 =  ( n296 ) ? ( n297 ) : ( n310 ) ;
assign n312 =  ( n294 ) ? ( n295 ) : ( n311 ) ;
assign n313 =  ( n291 ) ? ( n293 ) : ( n312 ) ;
assign n314 =  ( n304 ) ? ( n303 ) : ( n305 ) ;
assign n315 =  ( n302 ) ? ( n301 ) : ( n314 ) ;
assign n316 =  ( n300 ) ? ( n299 ) : ( n315 ) ;
assign n317 =  ( n298 ) ? ( n297 ) : ( n316 ) ;
assign n318 =  ( n296 ) ? ( n295 ) : ( n317 ) ;
assign n319 =  ( n294 ) ? ( n293 ) : ( n318 ) ;
assign n320 =  ( n291 ) ? ( n306 ) : ( n319 ) ;
assign n321 =  ( n304 ) ? ( n301 ) : ( n303 ) ;
assign n322 =  ( n302 ) ? ( n299 ) : ( n321 ) ;
assign n323 =  ( n300 ) ? ( n297 ) : ( n322 ) ;
assign n324 =  ( n298 ) ? ( n295 ) : ( n323 ) ;
assign n325 =  ( n296 ) ? ( n293 ) : ( n324 ) ;
assign n326 =  ( n294 ) ? ( n306 ) : ( n325 ) ;
assign n327 =  ( n291 ) ? ( n305 ) : ( n326 ) ;
assign n328 =  ( n304 ) ? ( n299 ) : ( n301 ) ;
assign n329 =  ( n302 ) ? ( n297 ) : ( n328 ) ;
assign n330 =  ( n300 ) ? ( n295 ) : ( n329 ) ;
assign n331 =  ( n298 ) ? ( n293 ) : ( n330 ) ;
assign n332 =  ( n296 ) ? ( n306 ) : ( n331 ) ;
assign n333 =  ( n294 ) ? ( n305 ) : ( n332 ) ;
assign n334 =  ( n291 ) ? ( n303 ) : ( n333 ) ;
assign n335 =  ( n304 ) ? ( n297 ) : ( n299 ) ;
assign n336 =  ( n302 ) ? ( n295 ) : ( n335 ) ;
assign n337 =  ( n300 ) ? ( n293 ) : ( n336 ) ;
assign n338 =  ( n298 ) ? ( n306 ) : ( n337 ) ;
assign n339 =  ( n296 ) ? ( n305 ) : ( n338 ) ;
assign n340 =  ( n294 ) ? ( n303 ) : ( n339 ) ;
assign n341 =  ( n291 ) ? ( n301 ) : ( n340 ) ;
assign n342 =  ( n304 ) ? ( n295 ) : ( n297 ) ;
assign n343 =  ( n302 ) ? ( n293 ) : ( n342 ) ;
assign n344 =  ( n300 ) ? ( n306 ) : ( n343 ) ;
assign n345 =  ( n298 ) ? ( n305 ) : ( n344 ) ;
assign n346 =  ( n296 ) ? ( n303 ) : ( n345 ) ;
assign n347 =  ( n294 ) ? ( n301 ) : ( n346 ) ;
assign n348 =  ( n291 ) ? ( n299 ) : ( n347 ) ;
assign n349 =  ( n304 ) ? ( n293 ) : ( n295 ) ;
assign n350 =  ( n302 ) ? ( n306 ) : ( n349 ) ;
assign n351 =  ( n300 ) ? ( n305 ) : ( n350 ) ;
assign n352 =  ( n298 ) ? ( n303 ) : ( n351 ) ;
assign n353 =  ( n296 ) ? ( n301 ) : ( n352 ) ;
assign n354 =  ( n294 ) ? ( n299 ) : ( n353 ) ;
assign n355 =  ( n291 ) ? ( n297 ) : ( n354 ) ;
assign n356 =  ( n304 ) ? ( n306 ) : ( n293 ) ;
assign n357 =  ( n302 ) ? ( n305 ) : ( n356 ) ;
assign n358 =  ( n300 ) ? ( n303 ) : ( n357 ) ;
assign n359 =  ( n298 ) ? ( n301 ) : ( n358 ) ;
assign n360 =  ( n296 ) ? ( n299 ) : ( n359 ) ;
assign n361 =  ( n294 ) ? ( n297 ) : ( n360 ) ;
assign n362 =  ( n291 ) ? ( n295 ) : ( n361 ) ;
assign n363 =  { ( n355 ) , ( n362 ) }  ;
assign n364 =  { ( n348 ) , ( n363 ) }  ;
assign n365 =  { ( n341 ) , ( n364 ) }  ;
assign n366 =  { ( n334 ) , ( n365 ) }  ;
assign n367 =  { ( n327 ) , ( n366 ) }  ;
assign n368 =  { ( n320 ) , ( n367 ) }  ;
assign n369 =  { ( n313 ) , ( n368 ) }  ;
assign n370 =  { ( pre_pix ) , ( n369 ) }  ;
assign n371 =  ( n232 ) ? ( stencil_8 ) : ( n370 ) ;
assign n372 =  ( n24 ) ? ( stencil_8 ) : ( stencil_8 ) ;
assign n373 =  ( n13 ) ? ( n371 ) : ( n372 ) ;
assign n374 =  ( n10 ) ? ( stencil_8 ) : ( n373 ) ;
assign n375 =  ( n4 ) ? ( stencil_8 ) : ( n374 ) ;
assign n376 = ~ ( n4 ) ;
assign n377 = ~ ( n10 ) ;
assign n378 =  ( n376 ) & ( n377 )  ;
assign n379 = ~ ( n13 ) ;
assign n380 =  ( n378 ) & ( n379 )  ;
assign n381 = ~ ( n24 ) ;
assign n382 =  ( n380 ) & ( n381 )  ;
assign n383 =  ( n380 ) & ( n24 )  ;
assign n384 =  ( n378 ) & ( n13 )  ;
assign n385 = ~ ( n291 ) ;
assign n386 =  ( n384 ) & ( n385 )  ;
assign n387 =  ( n384 ) & ( n291 )  ;
assign n388 =  ( n376 ) & ( n10 )  ;
assign RAM_0_addr0 = n387 ? (n292) : (0);
assign RAM_0_data0 = n387 ? (pre_pix) : (RAM_0[0]);
assign n389 = ~ ( n294 ) ;
assign n390 =  ( n384 ) & ( n389 )  ;
assign n391 =  ( n384 ) & ( n294 )  ;
assign RAM_1_addr0 = n391 ? (n292) : (0);
assign RAM_1_data0 = n391 ? (pre_pix) : (RAM_1[0]);
assign n392 = ~ ( n296 ) ;
assign n393 =  ( n384 ) & ( n392 )  ;
assign n394 =  ( n384 ) & ( n296 )  ;
assign RAM_2_addr0 = n394 ? (n292) : (0);
assign RAM_2_data0 = n394 ? (pre_pix) : (RAM_2[0]);
assign n395 = ~ ( n298 ) ;
assign n396 =  ( n384 ) & ( n395 )  ;
assign n397 =  ( n384 ) & ( n298 )  ;
assign RAM_3_addr0 = n397 ? (n292) : (0);
assign RAM_3_data0 = n397 ? (pre_pix) : (RAM_3[0]);
assign n398 = ~ ( n300 ) ;
assign n399 =  ( n384 ) & ( n398 )  ;
assign n400 =  ( n384 ) & ( n300 )  ;
assign RAM_4_addr0 = n400 ? (n292) : (0);
assign RAM_4_data0 = n400 ? (pre_pix) : (RAM_4[0]);
assign n401 = ~ ( n302 ) ;
assign n402 =  ( n384 ) & ( n401 )  ;
assign n403 =  ( n384 ) & ( n302 )  ;
assign RAM_5_addr0 = n403 ? (n292) : (0);
assign RAM_5_data0 = n403 ? (pre_pix) : (RAM_5[0]);
assign n404 = ~ ( n304 ) ;
assign n405 =  ( n384 ) & ( n404 )  ;
assign n406 =  ( n384 ) & ( n304 )  ;
assign RAM_6_addr0 = n406 ? (n292) : (0);
assign RAM_6_data0 = n406 ? (pre_pix) : (RAM_6[0]);
assign n407 = ~ ( n15 ) ;
assign n408 =  ( n384 ) & ( n407 )  ;
assign n409 =  ( n384 ) & ( n15 )  ;
assign RAM_7_addr0 = n409 ? (n292) : (0);
assign RAM_7_data0 = n409 ? (pre_pix) : (RAM_7[0]);
/*
function [7:0] gb_fun ;
input [647:0] arg0;
    begin
//TODO: Add the specific function HERE.    end
endfunction
*/

always @(posedge clk) begin
   if(rst) begin
       RAM_w <= RAM_w;
       RAM_x <= RAM_x;
       RAM_y <= RAM_y;
       arg_0_TDATA <= arg_0_TDATA;
       arg_0_TVALID <= arg_0_TVALID;
       arg_1_TREADY <= arg_1_TREADY;
       cur_pix <= cur_pix;
       gbit <= gbit;
       pre_pix <= pre_pix;
       proc_in <= proc_in;
       st_ready <= st_ready;
       stencil_0 <= stencil_0;
       stencil_1 <= stencil_1;
       stencil_2 <= stencil_2;
       stencil_3 <= stencil_3;
       stencil_4 <= stencil_4;
       stencil_5 <= stencil_5;
       stencil_6 <= stencil_6;
       stencil_7 <= stencil_7;
       stencil_8 <= stencil_8;
   end
   else if(step) begin
       RAM_w <= n28;
       RAM_x <= n34;
       RAM_y <= n42;
       arg_0_TDATA <= n219;
       arg_0_TVALID <= n225;
       arg_1_TREADY <= n237;
       cur_pix <= n241;
       gbit <= gbit;
       pre_pix <= n244;
       proc_in <= n247;
       st_ready <= n250;
       stencil_0 <= n255;
       stencil_1 <= n260;
       stencil_2 <= n265;
       stencil_3 <= n270;
       stencil_4 <= n275;
       stencil_5 <= n280;
       stencil_6 <= n285;
       stencil_7 <= n290;
       stencil_8 <= n375;
       RAM_0 [ RAM_0_addr0 ] <= RAM_0_data0;
       RAM_1 [ RAM_1_addr0 ] <= RAM_1_data0;
       RAM_2 [ RAM_2_addr0 ] <= RAM_2_data0;
       RAM_3 [ RAM_3_addr0 ] <= RAM_3_data0;
       RAM_4 [ RAM_4_addr0 ] <= RAM_4_data0;
       RAM_5 [ RAM_5_addr0 ] <= RAM_5_data0;
       RAM_6 [ RAM_6_addr0 ] <= RAM_6_data0;
       RAM_7 [ RAM_7_addr0 ] <= RAM_7_data0;
   end
end
endmodule
