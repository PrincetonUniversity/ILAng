module SPEC_B(
arg_0_TREADY,
arg_1_TDATA,
arg_1_TVALID,
LB1D_buff,
LB1D_in,
LB1D_it_1,
LB1D_p_cnt,
LB1D_uIn,
LB2D_proc_w,
LB2D_proc_x,
LB2D_proc_y,
LB2D_shift_0,
LB2D_shift_1,
LB2D_shift_2,
LB2D_shift_3,
LB2D_shift_4,
LB2D_shift_5,
LB2D_shift_6,
LB2D_shift_7,
LB2D_shift_x,
LB2D_shift_y,
arg_0_TDATA,
arg_0_TVALID,
arg_1_TREADY,
gb_exit_it_1,
gb_exit_it_2,
gb_exit_it_3,
gb_exit_it_4,
gb_exit_it_5,
gb_exit_it_6,
gb_exit_it_7,
gb_exit_it_8,
gb_p_cnt,
gb_pp_it_1,
gb_pp_it_2,
gb_pp_it_3,
gb_pp_it_4,
gb_pp_it_5,
gb_pp_it_6,
gb_pp_it_7,
gb_pp_it_8,
gb_pp_it_9,
in_stream_buff_0,
in_stream_buff_1,
in_stream_empty,
in_stream_full,
slice_stream_buff_0,
slice_stream_buff_1,
slice_stream_empty,
slice_stream_full,
stencil_stream_buff_0,
stencil_stream_buff_1,
stencil_stream_empty,
stencil_stream_full,
clk,rst,
step
);
input            arg_0_TREADY;
input      [7:0] arg_1_TDATA;
input            arg_1_TVALID;
input clk;
input rst;
input step;
output      [7:0] LB1D_buff;
output      [7:0] LB1D_in;
output            LB1D_it_1;
output     [18:0] LB1D_p_cnt;
output      [7:0] LB1D_uIn;
output     [63:0] LB2D_proc_w;
output      [8:0] LB2D_proc_x;
output      [9:0] LB2D_proc_y;
output     [71:0] LB2D_shift_0;
output     [71:0] LB2D_shift_1;
output     [71:0] LB2D_shift_2;
output     [71:0] LB2D_shift_3;
output     [71:0] LB2D_shift_4;
output     [71:0] LB2D_shift_5;
output     [71:0] LB2D_shift_6;
output     [71:0] LB2D_shift_7;
output      [8:0] LB2D_shift_x;
output      [9:0] LB2D_shift_y;
output      [7:0] arg_0_TDATA;
output            arg_0_TVALID;
output            arg_1_TREADY;
output            gb_exit_it_1;
output            gb_exit_it_2;
output            gb_exit_it_3;
output            gb_exit_it_4;
output            gb_exit_it_5;
output            gb_exit_it_6;
output            gb_exit_it_7;
output            gb_exit_it_8;
output     [18:0] gb_p_cnt;
output            gb_pp_it_1;
output            gb_pp_it_2;
output            gb_pp_it_3;
output            gb_pp_it_4;
output            gb_pp_it_5;
output            gb_pp_it_6;
output            gb_pp_it_7;
output            gb_pp_it_8;
output            gb_pp_it_9;
output      [7:0] in_stream_buff_0;
output      [7:0] in_stream_buff_1;
output            in_stream_empty;
output            in_stream_full;
output     [71:0] slice_stream_buff_0;
output     [71:0] slice_stream_buff_1;
output            slice_stream_empty;
output            slice_stream_full;
output    [647:0] stencil_stream_buff_0;
output    [647:0] stencil_stream_buff_1;
output            stencil_stream_empty;
output            stencil_stream_full;
reg      [7:0] LB1D_buff;
reg      [7:0] LB1D_in;
reg            LB1D_it_1;
reg     [18:0] LB1D_p_cnt;
reg      [7:0] LB1D_uIn;
reg     [63:0] LB2D_proc_w;
reg      [8:0] LB2D_proc_x;
reg      [9:0] LB2D_proc_y;
reg     [71:0] LB2D_shift_0;
reg     [71:0] LB2D_shift_1;
reg     [71:0] LB2D_shift_2;
reg     [71:0] LB2D_shift_3;
reg     [71:0] LB2D_shift_4;
reg     [71:0] LB2D_shift_5;
reg     [71:0] LB2D_shift_6;
reg     [71:0] LB2D_shift_7;
reg      [8:0] LB2D_shift_x;
reg      [9:0] LB2D_shift_y;
reg      [7:0] arg_0_TDATA;
reg            arg_0_TVALID;
reg            arg_1_TREADY;
reg            gb_exit_it_1;
reg            gb_exit_it_2;
reg            gb_exit_it_3;
reg            gb_exit_it_4;
reg            gb_exit_it_5;
reg            gb_exit_it_6;
reg            gb_exit_it_7;
reg            gb_exit_it_8;
reg     [18:0] gb_p_cnt;
reg            gb_pp_it_1;
reg            gb_pp_it_2;
reg            gb_pp_it_3;
reg            gb_pp_it_4;
reg            gb_pp_it_5;
reg            gb_pp_it_6;
reg            gb_pp_it_7;
reg            gb_pp_it_8;
reg            gb_pp_it_9;
reg      [7:0] in_stream_buff_0;
reg      [7:0] in_stream_buff_1;
reg            in_stream_empty;
reg            in_stream_full;
reg     [71:0] slice_stream_buff_0;
reg     [71:0] slice_stream_buff_1;
reg            slice_stream_empty;
reg            slice_stream_full;
reg    [647:0] stencil_stream_buff_0;
reg    [647:0] stencil_stream_buff_1;
reg            stencil_stream_empty;
reg            stencil_stream_full;
wire            arg_0_TREADY;
wire      [7:0] arg_1_TDATA;
wire            arg_1_TVALID;
wire            n0;
wire            n1;
wire            n2;
wire            n3;
wire            n4;
wire            n5;
wire            n6;
wire            n7;
wire            n8;
wire            n9;
wire            n10;
wire            n11;
wire            n12;
wire            n13;
wire            n14;
wire            n15;
wire            n16;
wire            n17;
wire            n18;
wire            n19;
wire            n20;
wire            n21;
wire            n22;
wire            n23;
wire            n24;
wire            n25;
wire            n26;
wire            n27;
wire            n28;
wire            n29;
wire            n30;
wire            n31;
wire            n32;
wire            n33;
wire            n34;
wire            n35;
wire            n36;
wire            n37;
wire            n38;
wire            n39;
wire      [7:0] n40;
wire      [7:0] n41;
wire      [7:0] n42;
wire      [7:0] n43;
wire      [7:0] n44;
wire      [7:0] n45;
wire      [7:0] n46;
wire      [7:0] n47;
wire      [7:0] n48;
wire      [7:0] n49;
wire      [7:0] n50;
wire      [7:0] n51;
wire      [7:0] n52;
wire      [7:0] n53;
wire            n54;
wire            n55;
wire            n56;
wire     [18:0] n57;
wire     [18:0] n58;
wire     [18:0] n59;
wire     [18:0] n60;
wire     [18:0] n61;
wire     [18:0] n62;
wire     [18:0] n63;
wire     [18:0] n64;
wire      [7:0] n65;
wire      [7:0] n66;
wire      [7:0] n67;
wire      [7:0] n68;
wire      [7:0] n69;
wire      [7:0] n70;
wire            n71;
wire            n72;
wire     [63:0] n73;
wire     [63:0] n74;
wire     [63:0] n75;
wire     [63:0] n76;
wire     [63:0] n77;
wire     [63:0] n78;
wire     [63:0] n79;
wire     [63:0] n80;
wire     [63:0] n81;
wire      [8:0] n82;
wire      [8:0] n83;
wire      [8:0] n84;
wire      [8:0] n85;
wire      [8:0] n86;
wire      [8:0] n87;
wire      [8:0] n88;
wire      [8:0] n89;
wire            n90;
wire      [9:0] n91;
wire      [9:0] n92;
wire      [9:0] n93;
wire      [9:0] n94;
wire      [9:0] n95;
wire      [9:0] n96;
wire      [9:0] n97;
wire      [9:0] n98;
wire      [9:0] n99;
wire     [71:0] n100;
wire     [71:0] n101;
wire     [71:0] n102;
wire     [71:0] n103;
wire     [71:0] n104;
wire     [71:0] n105;
wire     [71:0] n106;
wire     [71:0] n107;
wire     [71:0] n108;
wire     [71:0] n109;
wire     [71:0] n110;
wire     [71:0] n111;
wire     [71:0] n112;
wire     [71:0] n113;
wire     [71:0] n114;
wire     [71:0] n115;
wire     [71:0] n116;
wire     [71:0] n117;
wire     [71:0] n118;
wire     [71:0] n119;
wire     [71:0] n120;
wire     [71:0] n121;
wire     [71:0] n122;
wire     [71:0] n123;
wire     [71:0] n124;
wire     [71:0] n125;
wire     [71:0] n126;
wire     [71:0] n127;
wire     [71:0] n128;
wire     [71:0] n129;
wire     [71:0] n130;
wire     [71:0] n131;
wire     [71:0] n132;
wire     [71:0] n133;
wire     [71:0] n134;
wire     [71:0] n135;
wire     [71:0] n136;
wire     [71:0] n137;
wire     [71:0] n138;
wire     [71:0] n139;
wire     [71:0] n140;
wire     [71:0] n141;
wire            n142;
wire     [71:0] n143;
wire     [71:0] n144;
wire     [71:0] n145;
wire     [71:0] n146;
wire     [71:0] n147;
wire     [71:0] n148;
wire     [71:0] n149;
wire            n150;
wire            n151;
wire            n152;
wire            n153;
wire      [8:0] n154;
wire      [8:0] n155;
wire      [8:0] n156;
wire      [8:0] n157;
wire      [8:0] n158;
wire      [8:0] n159;
wire      [8:0] n160;
wire      [8:0] n161;
wire            n162;
wire            n163;
wire      [9:0] n164;
wire      [9:0] n165;
wire      [9:0] n166;
wire      [9:0] n167;
wire      [9:0] n168;
wire      [9:0] n169;
wire      [9:0] n170;
wire      [9:0] n171;
wire      [9:0] n172;
wire            n173;
wire    [647:0] n174;
wire      [7:0] n175;
wire      [7:0] n176;
wire      [7:0] n177;
wire      [7:0] n178;
wire      [7:0] n179;
wire      [7:0] n180;
wire      [7:0] n181;
wire            n182;
wire            n183;
wire            n184;
wire            n185;
wire            n186;
wire            n187;
wire            n188;
wire            n189;
wire            n190;
wire            n191;
wire            n192;
wire            n193;
wire            n194;
wire            n195;
wire            n196;
wire            n197;
wire            n198;
wire            n199;
wire            n200;
wire            n201;
wire            n202;
wire            n203;
wire            n204;
wire            n205;
wire            n206;
wire            n207;
wire            n208;
wire            n209;
wire            n210;
wire            n211;
wire            n212;
wire            n213;
wire            n214;
wire            n215;
wire            n216;
wire            n217;
wire            n218;
wire            n219;
wire            n220;
wire            n221;
wire            n222;
wire            n223;
wire            n224;
wire            n225;
wire            n226;
wire            n227;
wire            n228;
wire            n229;
wire            n230;
wire            n231;
wire            n232;
wire            n233;
wire            n234;
wire            n235;
wire            n236;
wire            n237;
wire            n238;
wire            n239;
wire            n240;
wire            n241;
wire            n242;
wire            n243;
wire            n244;
wire            n245;
wire            n246;
wire            n247;
wire            n248;
wire     [18:0] n249;
wire     [18:0] n250;
wire     [18:0] n251;
wire     [18:0] n252;
wire     [18:0] n253;
wire     [18:0] n254;
wire     [18:0] n255;
wire     [18:0] n256;
wire            n257;
wire            n258;
wire            n259;
wire            n260;
wire            n261;
wire            n262;
wire            n263;
wire            n264;
wire            n265;
wire            n266;
wire            n267;
wire            n268;
wire            n269;
wire            n270;
wire            n271;
wire            n272;
wire            n273;
wire            n274;
wire            n275;
wire            n276;
wire            n277;
wire            n278;
wire            n279;
wire            n280;
wire            n281;
wire            n282;
wire            n283;
wire            n284;
wire            n285;
wire            n286;
wire            n287;
wire            n288;
wire            n289;
wire            n290;
wire            n291;
wire            n292;
wire            n293;
wire            n294;
wire            n295;
wire            n296;
wire            n297;
wire            n298;
wire            n299;
wire            n300;
wire            n301;
wire            n302;
wire            n303;
wire            n304;
wire            n305;
wire            n306;
wire            n307;
wire            n308;
wire            n309;
wire            n310;
wire      [7:0] n311;
wire      [7:0] n312;
wire      [7:0] n313;
wire      [7:0] n314;
wire      [7:0] n315;
wire      [7:0] n316;
wire      [7:0] n317;
wire      [7:0] n318;
wire      [7:0] n319;
wire      [7:0] n320;
wire      [7:0] n321;
wire      [7:0] n322;
wire            n323;
wire            n324;
wire            n325;
wire            n326;
wire            n327;
wire            n328;
wire            n329;
wire            n330;
wire            n331;
wire            n332;
wire            n333;
wire            n334;
wire            n335;
wire            n336;
wire            n337;
wire            n338;
wire      [7:0] n339;
wire            n340;
wire      [8:0] n341;
wire      [7:0] n342;
wire            n343;
wire      [7:0] n344;
wire            n345;
wire      [7:0] n346;
wire            n347;
wire      [7:0] n348;
wire            n349;
wire      [7:0] n350;
wire            n351;
wire      [7:0] n352;
wire            n353;
wire      [7:0] n354;
wire      [7:0] n355;
wire      [7:0] n356;
wire      [7:0] n357;
wire      [7:0] n358;
wire      [7:0] n359;
wire      [7:0] n360;
wire      [7:0] n361;
wire      [7:0] n362;
wire      [7:0] n363;
wire      [7:0] n364;
wire      [7:0] n365;
wire      [7:0] n366;
wire      [7:0] n367;
wire      [7:0] n368;
wire      [7:0] n369;
wire      [7:0] n370;
wire      [7:0] n371;
wire      [7:0] n372;
wire      [7:0] n373;
wire      [7:0] n374;
wire      [7:0] n375;
wire      [7:0] n376;
wire      [7:0] n377;
wire      [7:0] n378;
wire      [7:0] n379;
wire      [7:0] n380;
wire      [7:0] n381;
wire      [7:0] n382;
wire      [7:0] n383;
wire      [7:0] n384;
wire      [7:0] n385;
wire      [7:0] n386;
wire      [7:0] n387;
wire      [7:0] n388;
wire      [7:0] n389;
wire      [7:0] n390;
wire      [7:0] n391;
wire      [7:0] n392;
wire      [7:0] n393;
wire      [7:0] n394;
wire      [7:0] n395;
wire      [7:0] n396;
wire      [7:0] n397;
wire      [7:0] n398;
wire      [7:0] n399;
wire      [7:0] n400;
wire      [7:0] n401;
wire      [7:0] n402;
wire      [7:0] n403;
wire      [7:0] n404;
wire      [7:0] n405;
wire      [7:0] n406;
wire      [7:0] n407;
wire      [7:0] n408;
wire      [7:0] n409;
wire      [7:0] n410;
wire      [7:0] n411;
wire     [15:0] n412;
wire     [23:0] n413;
wire     [31:0] n414;
wire     [39:0] n415;
wire     [47:0] n416;
wire     [55:0] n417;
wire     [63:0] n418;
wire     [71:0] n419;
wire     [71:0] n420;
wire     [71:0] n421;
wire     [71:0] n422;
wire     [71:0] n423;
wire     [71:0] n424;
wire     [71:0] n425;
wire     [71:0] n426;
wire     [71:0] n427;
wire     [71:0] n428;
wire     [71:0] n429;
wire     [71:0] n430;
wire     [71:0] n431;
wire     [71:0] n432;
wire     [71:0] n433;
wire            n434;
wire            n435;
wire            n436;
wire            n437;
wire            n438;
wire            n439;
wire            n440;
wire            n441;
wire            n442;
wire            n443;
wire            n444;
wire            n445;
wire            n446;
wire            n447;
wire            n448;
wire            n449;
wire            n450;
wire            n451;
wire            n452;
wire            n453;
wire      [7:0] n454;
wire      [7:0] n455;
wire      [7:0] n456;
wire      [7:0] n457;
wire      [7:0] n458;
wire      [7:0] n459;
wire      [7:0] n460;
wire      [7:0] n461;
wire      [7:0] n462;
wire     [15:0] n463;
wire     [23:0] n464;
wire     [31:0] n465;
wire     [39:0] n466;
wire     [47:0] n467;
wire     [55:0] n468;
wire     [63:0] n469;
wire     [71:0] n470;
wire      [7:0] n471;
wire      [7:0] n472;
wire      [7:0] n473;
wire      [7:0] n474;
wire      [7:0] n475;
wire      [7:0] n476;
wire      [7:0] n477;
wire      [7:0] n478;
wire      [7:0] n479;
wire     [15:0] n480;
wire     [23:0] n481;
wire     [31:0] n482;
wire     [39:0] n483;
wire     [47:0] n484;
wire     [55:0] n485;
wire     [63:0] n486;
wire     [71:0] n487;
wire      [7:0] n488;
wire      [7:0] n489;
wire      [7:0] n490;
wire      [7:0] n491;
wire      [7:0] n492;
wire      [7:0] n493;
wire      [7:0] n494;
wire      [7:0] n495;
wire      [7:0] n496;
wire     [15:0] n497;
wire     [23:0] n498;
wire     [31:0] n499;
wire     [39:0] n500;
wire     [47:0] n501;
wire     [55:0] n502;
wire     [63:0] n503;
wire     [71:0] n504;
wire      [7:0] n505;
wire      [7:0] n506;
wire      [7:0] n507;
wire      [7:0] n508;
wire      [7:0] n509;
wire      [7:0] n510;
wire      [7:0] n511;
wire      [7:0] n512;
wire      [7:0] n513;
wire     [15:0] n514;
wire     [23:0] n515;
wire     [31:0] n516;
wire     [39:0] n517;
wire     [47:0] n518;
wire     [55:0] n519;
wire     [63:0] n520;
wire     [71:0] n521;
wire      [7:0] n522;
wire      [7:0] n523;
wire      [7:0] n524;
wire      [7:0] n525;
wire      [7:0] n526;
wire      [7:0] n527;
wire      [7:0] n528;
wire      [7:0] n529;
wire      [7:0] n530;
wire     [15:0] n531;
wire     [23:0] n532;
wire     [31:0] n533;
wire     [39:0] n534;
wire     [47:0] n535;
wire     [55:0] n536;
wire     [63:0] n537;
wire     [71:0] n538;
wire      [7:0] n539;
wire      [7:0] n540;
wire      [7:0] n541;
wire      [7:0] n542;
wire      [7:0] n543;
wire      [7:0] n544;
wire      [7:0] n545;
wire      [7:0] n546;
wire      [7:0] n547;
wire     [15:0] n548;
wire     [23:0] n549;
wire     [31:0] n550;
wire     [39:0] n551;
wire     [47:0] n552;
wire     [55:0] n553;
wire     [63:0] n554;
wire     [71:0] n555;
wire      [7:0] n556;
wire      [7:0] n557;
wire      [7:0] n558;
wire      [7:0] n559;
wire      [7:0] n560;
wire      [7:0] n561;
wire      [7:0] n562;
wire      [7:0] n563;
wire      [7:0] n564;
wire     [15:0] n565;
wire     [23:0] n566;
wire     [31:0] n567;
wire     [39:0] n568;
wire     [47:0] n569;
wire     [55:0] n570;
wire     [63:0] n571;
wire     [71:0] n572;
wire      [7:0] n573;
wire      [7:0] n574;
wire      [7:0] n575;
wire      [7:0] n576;
wire      [7:0] n577;
wire      [7:0] n578;
wire      [7:0] n579;
wire      [7:0] n580;
wire      [7:0] n581;
wire     [15:0] n582;
wire     [23:0] n583;
wire     [31:0] n584;
wire     [39:0] n585;
wire     [47:0] n586;
wire     [55:0] n587;
wire     [63:0] n588;
wire     [71:0] n589;
wire      [7:0] n590;
wire      [7:0] n591;
wire      [7:0] n592;
wire      [7:0] n593;
wire      [7:0] n594;
wire      [7:0] n595;
wire      [7:0] n596;
wire      [7:0] n597;
wire      [7:0] n598;
wire     [15:0] n599;
wire     [23:0] n600;
wire     [31:0] n601;
wire     [39:0] n602;
wire     [47:0] n603;
wire     [55:0] n604;
wire     [63:0] n605;
wire     [71:0] n606;
wire    [143:0] n607;
wire    [215:0] n608;
wire    [287:0] n609;
wire    [359:0] n610;
wire    [431:0] n611;
wire    [503:0] n612;
wire    [575:0] n613;
wire    [647:0] n614;
wire    [647:0] n615;
wire    [647:0] n616;
wire    [647:0] n617;
wire    [647:0] n618;
wire    [647:0] n619;
wire    [647:0] n620;
wire    [647:0] n621;
wire    [647:0] n622;
wire    [647:0] n623;
wire    [647:0] n624;
wire    [647:0] n625;
wire    [647:0] n626;
wire    [647:0] n627;
wire            n628;
wire            n629;
wire            n630;
wire            n631;
wire            n632;
wire            n633;
wire            n634;
wire            n635;
wire            n636;
wire            n637;
wire            n638;
wire            n639;
wire            n640;
wire            n641;
wire            n642;
wire            n643;
wire            n644;
wire            n645;
wire            n646;
wire      [8:0] LB2D_proc_0_addr0;
wire      [7:0] LB2D_proc_0_data0;
wire            n647;
wire            n648;
wire            n649;
wire            n650;
wire            n651;
wire            n652;
wire            n653;
wire            n654;
wire            n655;
wire            n656;
wire            n657;
wire            n658;
wire            n659;
wire            n660;
wire            n661;
wire            n662;
wire            n663;
wire            n664;
wire            n665;
wire      [8:0] LB2D_proc_1_addr0;
wire      [7:0] LB2D_proc_1_data0;
wire            n666;
wire            n667;
wire            n668;
wire      [8:0] LB2D_proc_2_addr0;
wire      [7:0] LB2D_proc_2_data0;
wire            n669;
wire            n670;
wire            n671;
wire      [8:0] LB2D_proc_3_addr0;
wire      [7:0] LB2D_proc_3_data0;
wire            n672;
wire            n673;
wire            n674;
wire      [8:0] LB2D_proc_4_addr0;
wire      [7:0] LB2D_proc_4_data0;
wire            n675;
wire            n676;
wire            n677;
wire      [8:0] LB2D_proc_5_addr0;
wire      [7:0] LB2D_proc_5_data0;
wire            n678;
wire            n679;
wire            n680;
wire      [8:0] LB2D_proc_6_addr0;
wire      [7:0] LB2D_proc_6_data0;
wire            n681;
wire            n682;
wire            n683;
wire      [8:0] LB2D_proc_7_addr0;
wire      [7:0] LB2D_proc_7_data0;
wire            n684;
wire            n685;
wire            n686;
reg      [7:0] LB2D_proc_0[511:0];
reg      [7:0] LB2D_proc_1[511:0];
reg      [7:0] LB2D_proc_2[511:0];
reg      [7:0] LB2D_proc_3[511:0];
reg      [7:0] LB2D_proc_4[511:0];
reg      [7:0] LB2D_proc_5[511:0];
reg      [7:0] LB2D_proc_6[511:0];
reg      [7:0] LB2D_proc_7[511:0];
wire clk;
wire rst;
wire step;
assign n0 =  ( arg_1_TREADY ) == ( 1'd1 )  ;
assign n1 =  ( in_stream_full ) == ( 1'd0 )  ;
assign n2 =  ( n0 ) & ( n1 )  ;
assign n3 =  ( LB1D_it_1 ) == ( 1'd1 )  ;
assign n4 =  ( n2 ) & ( n3 )  ;
assign n5 =  ( LB1D_p_cnt ) == ( 19'd316224 )  ;
assign n6 =  ( n4 ) & ( n5 )  ;
assign n7 =  ( arg_0_TREADY ) == ( 1'd1 )  ;
assign n8 =  ( arg_0_TVALID ) == ( 1'd1 )  ;
assign n9 =  ( n7 ) & ( n8 )  ;
assign n10 =  ( arg_1_TVALID ) == ( 1'd0 )  ;
assign n11 =  ( n9 ) & ( n10 )  ;
assign n12 =  ( arg_0_TVALID ) == ( 1'd0 )  ;
assign n13 =  ( gb_exit_it_1 ) == ( 1'd0 )  ;
assign n14 =  ( stencil_stream_empty ) == ( 1'd0 )  ;
assign n15 =  ( n13 ) & ( n14 )  ;
assign n16 =  ( gb_exit_it_1 ) == ( 1'd1 )  ;
assign n17 =  ( gb_exit_it_8 ) == ( 1'd0 )  ;
assign n18 =  ( n16 ) & ( n17 )  ;
assign n19 =  ( n15 ) | ( n18 )  ;
assign n20 =  ( n12 ) & ( n19 )  ;
assign n21 =  ( slice_stream_empty ) == ( 1'd0 )  ;
assign n22 =  ( LB2D_shift_x ) != ( 9'd488 )  ;
assign n23 =  ( n21 ) & ( n22 )  ;
assign n24 =  ( stencil_stream_full ) == ( 1'd0 )  ;
assign n25 =  ( LB2D_shift_x ) < ( 9'd8 )  ;
assign n26 =  ( LB2D_shift_x ) > ( 9'd0 )  ;
assign n27 =  ( n25 ) & ( n26 )  ;
assign n28 =  ( n24 ) | ( n27 )  ;
assign n29 =  ( n23 ) & ( n28 )  ;
assign n30 =  ( in_stream_empty ) == ( 1'd0 )  ;
assign n31 =  ( slice_stream_full ) == ( 1'd0 )  ;
assign n32 =  ( LB2D_proc_y ) < ( 10'd8 )  ;
assign n33 =  ( n31 ) | ( n32 )  ;
assign n34 =  ( n30 ) & ( n33 )  ;
assign n35 =  ( arg_1_TREADY ) == ( 1'd0 )  ;
assign n36 =  ( n35 ) & ( n1 )  ;
assign n37 =  ( LB1D_it_1 ) == ( 1'd0 )  ;
assign n38 =  ( n36 ) & ( n37 )  ;
assign n39 =  ( n36 ) & ( n3 )  ;
assign n40 =  ( n39 ) ? ( LB1D_uIn ) : ( LB1D_buff ) ;
assign n41 =  ( n38 ) ? ( LB1D_uIn ) : ( n40 ) ;
assign n42 =  ( n34 ) ? ( LB1D_buff ) : ( n41 ) ;
assign n43 =  ( n29 ) ? ( LB1D_buff ) : ( n42 ) ;
assign n44 =  ( n20 ) ? ( LB1D_buff ) : ( n43 ) ;
assign n45 =  ( n11 ) ? ( LB1D_buff ) : ( n44 ) ;
assign n46 =  ( n6 ) ? ( LB1D_uIn ) : ( n45 ) ;
assign n47 =  ( n39 ) ? ( LB1D_in ) : ( LB1D_in ) ;
assign n48 =  ( n38 ) ? ( LB1D_in ) : ( n47 ) ;
assign n49 =  ( n34 ) ? ( LB1D_in ) : ( n48 ) ;
assign n50 =  ( n29 ) ? ( LB1D_in ) : ( n49 ) ;
assign n51 =  ( n20 ) ? ( LB1D_in ) : ( n50 ) ;
assign n52 =  ( n11 ) ? ( LB1D_in ) : ( n51 ) ;
assign n53 =  ( n6 ) ? ( LB1D_in ) : ( n52 ) ;
assign n54 =  ( n39 ) ? ( 1'd1 ) : ( LB1D_it_1 ) ;
assign n55 =  ( n38 ) ? ( 1'd1 ) : ( n54 ) ;
assign n56 =  ( n6 ) ? ( 1'd0 ) : ( n55 ) ;
assign n57 =  ( LB1D_p_cnt ) + ( 19'd1 )  ;
assign n58 =  ( n39 ) ? ( n57 ) : ( LB1D_p_cnt ) ;
assign n59 =  ( n38 ) ? ( n57 ) : ( n58 ) ;
assign n60 =  ( n34 ) ? ( LB1D_p_cnt ) : ( n59 ) ;
assign n61 =  ( n29 ) ? ( LB1D_p_cnt ) : ( n60 ) ;
assign n62 =  ( n20 ) ? ( LB1D_p_cnt ) : ( n61 ) ;
assign n63 =  ( n11 ) ? ( LB1D_p_cnt ) : ( n62 ) ;
assign n64 =  ( n6 ) ? ( 19'd0 ) : ( n63 ) ;
assign n65 =  ( n39 ) ? ( LB1D_in ) : ( LB1D_uIn ) ;
assign n66 =  ( n38 ) ? ( LB1D_in ) : ( n65 ) ;
assign n67 =  ( n34 ) ? ( LB1D_uIn ) : ( n66 ) ;
assign n68 =  ( n29 ) ? ( LB1D_uIn ) : ( n67 ) ;
assign n69 =  ( n20 ) ? ( LB1D_uIn ) : ( n68 ) ;
assign n70 =  ( n6 ) ? ( LB1D_in ) : ( n69 ) ;
assign n71 =  ( LB2D_proc_x ) == ( 9'd488 )  ;
assign n72 =  ( LB2D_proc_w ) == ( 64'd7 )  ;
assign n73 =  ( LB2D_proc_w ) + ( 64'd1 )  ;
assign n74 =  ( n72 ) ? ( 64'd0 ) : ( n73 ) ;
assign n75 =  ( n71 ) ? ( n74 ) : ( LB2D_proc_w ) ;
assign n76 =  ( n39 ) ? ( LB2D_proc_w ) : ( LB2D_proc_w ) ;
assign n77 =  ( n34 ) ? ( n75 ) : ( n76 ) ;
assign n78 =  ( n29 ) ? ( LB2D_proc_w ) : ( n77 ) ;
assign n79 =  ( n20 ) ? ( LB2D_proc_w ) : ( n78 ) ;
assign n80 =  ( n11 ) ? ( LB2D_proc_w ) : ( n79 ) ;
assign n81 =  ( n6 ) ? ( LB2D_proc_w ) : ( n80 ) ;
assign n82 =  ( LB2D_proc_x ) + ( 9'd1 )  ;
assign n83 =  ( n71 ) ? ( 9'd1 ) : ( n82 ) ;
assign n84 =  ( n39 ) ? ( LB2D_proc_x ) : ( LB2D_proc_x ) ;
assign n85 =  ( n34 ) ? ( n83 ) : ( n84 ) ;
assign n86 =  ( n29 ) ? ( LB2D_proc_x ) : ( n85 ) ;
assign n87 =  ( n20 ) ? ( LB2D_proc_x ) : ( n86 ) ;
assign n88 =  ( n11 ) ? ( LB2D_proc_x ) : ( n87 ) ;
assign n89 =  ( n6 ) ? ( LB2D_proc_x ) : ( n88 ) ;
assign n90 =  ( LB2D_proc_y ) == ( 10'd648 )  ;
assign n91 =  ( LB2D_proc_y ) + ( 10'd1 )  ;
assign n92 =  ( n90 ) ? ( 10'd0 ) : ( n91 ) ;
assign n93 =  ( n71 ) ? ( n92 ) : ( LB2D_proc_y ) ;
assign n94 =  ( n39 ) ? ( LB2D_proc_y ) : ( LB2D_proc_y ) ;
assign n95 =  ( n34 ) ? ( n93 ) : ( n94 ) ;
assign n96 =  ( n29 ) ? ( LB2D_proc_y ) : ( n95 ) ;
assign n97 =  ( n20 ) ? ( LB2D_proc_y ) : ( n96 ) ;
assign n98 =  ( n11 ) ? ( LB2D_proc_y ) : ( n97 ) ;
assign n99 =  ( n6 ) ? ( LB2D_proc_y ) : ( n98 ) ;
assign n100 =  ( n39 ) ? ( LB2D_shift_0 ) : ( LB2D_shift_0 ) ;
assign n101 =  ( n34 ) ? ( LB2D_shift_0 ) : ( n100 ) ;
assign n102 =  ( n29 ) ? ( LB2D_shift_1 ) : ( n101 ) ;
assign n103 =  ( n20 ) ? ( LB2D_shift_0 ) : ( n102 ) ;
assign n104 =  ( n11 ) ? ( LB2D_shift_0 ) : ( n103 ) ;
assign n105 =  ( n6 ) ? ( LB2D_shift_0 ) : ( n104 ) ;
assign n106 =  ( n39 ) ? ( LB2D_shift_1 ) : ( LB2D_shift_1 ) ;
assign n107 =  ( n34 ) ? ( LB2D_shift_1 ) : ( n106 ) ;
assign n108 =  ( n29 ) ? ( LB2D_shift_2 ) : ( n107 ) ;
assign n109 =  ( n20 ) ? ( LB2D_shift_1 ) : ( n108 ) ;
assign n110 =  ( n11 ) ? ( LB2D_shift_1 ) : ( n109 ) ;
assign n111 =  ( n6 ) ? ( LB2D_shift_1 ) : ( n110 ) ;
assign n112 =  ( n39 ) ? ( LB2D_shift_2 ) : ( LB2D_shift_2 ) ;
assign n113 =  ( n34 ) ? ( LB2D_shift_2 ) : ( n112 ) ;
assign n114 =  ( n29 ) ? ( LB2D_shift_3 ) : ( n113 ) ;
assign n115 =  ( n20 ) ? ( LB2D_shift_2 ) : ( n114 ) ;
assign n116 =  ( n11 ) ? ( LB2D_shift_2 ) : ( n115 ) ;
assign n117 =  ( n6 ) ? ( LB2D_shift_2 ) : ( n116 ) ;
assign n118 =  ( n39 ) ? ( LB2D_shift_3 ) : ( LB2D_shift_3 ) ;
assign n119 =  ( n34 ) ? ( LB2D_shift_3 ) : ( n118 ) ;
assign n120 =  ( n29 ) ? ( LB2D_shift_4 ) : ( n119 ) ;
assign n121 =  ( n20 ) ? ( LB2D_shift_3 ) : ( n120 ) ;
assign n122 =  ( n11 ) ? ( LB2D_shift_3 ) : ( n121 ) ;
assign n123 =  ( n6 ) ? ( LB2D_shift_3 ) : ( n122 ) ;
assign n124 =  ( n39 ) ? ( LB2D_shift_4 ) : ( LB2D_shift_4 ) ;
assign n125 =  ( n34 ) ? ( LB2D_shift_4 ) : ( n124 ) ;
assign n126 =  ( n29 ) ? ( LB2D_shift_5 ) : ( n125 ) ;
assign n127 =  ( n20 ) ? ( LB2D_shift_4 ) : ( n126 ) ;
assign n128 =  ( n11 ) ? ( LB2D_shift_4 ) : ( n127 ) ;
assign n129 =  ( n6 ) ? ( LB2D_shift_4 ) : ( n128 ) ;
assign n130 =  ( n39 ) ? ( LB2D_shift_5 ) : ( LB2D_shift_5 ) ;
assign n131 =  ( n34 ) ? ( LB2D_shift_5 ) : ( n130 ) ;
assign n132 =  ( n29 ) ? ( LB2D_shift_6 ) : ( n131 ) ;
assign n133 =  ( n20 ) ? ( LB2D_shift_5 ) : ( n132 ) ;
assign n134 =  ( n11 ) ? ( LB2D_shift_5 ) : ( n133 ) ;
assign n135 =  ( n6 ) ? ( LB2D_shift_5 ) : ( n134 ) ;
assign n136 =  ( n39 ) ? ( LB2D_shift_6 ) : ( LB2D_shift_6 ) ;
assign n137 =  ( n34 ) ? ( LB2D_shift_6 ) : ( n136 ) ;
assign n138 =  ( n29 ) ? ( LB2D_shift_7 ) : ( n137 ) ;
assign n139 =  ( n20 ) ? ( LB2D_shift_6 ) : ( n138 ) ;
assign n140 =  ( n11 ) ? ( LB2D_shift_6 ) : ( n139 ) ;
assign n141 =  ( n6 ) ? ( LB2D_shift_6 ) : ( n140 ) ;
assign n142 =  ( slice_stream_full ) == ( 1'd1 )  ;
assign n143 =  ( n142 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n144 =  ( n39 ) ? ( LB2D_shift_7 ) : ( LB2D_shift_7 ) ;
assign n145 =  ( n34 ) ? ( LB2D_shift_7 ) : ( n144 ) ;
assign n146 =  ( n29 ) ? ( n143 ) : ( n145 ) ;
assign n147 =  ( n20 ) ? ( LB2D_shift_7 ) : ( n146 ) ;
assign n148 =  ( n11 ) ? ( LB2D_shift_7 ) : ( n147 ) ;
assign n149 =  ( n6 ) ? ( LB2D_shift_7 ) : ( n148 ) ;
assign n150 =  ( LB2D_shift_x ) == ( 9'd488 )  ;
assign n151 =  ( n21 ) & ( n150 )  ;
assign n152 =  ( n24 ) | ( n25 )  ;
assign n153 =  ( n151 ) & ( n152 )  ;
assign n154 =  ( LB2D_shift_x ) + ( 9'd1 )  ;
assign n155 =  ( n39 ) ? ( LB2D_shift_x ) : ( LB2D_shift_x ) ;
assign n156 =  ( n34 ) ? ( LB2D_shift_x ) : ( n155 ) ;
assign n157 =  ( n29 ) ? ( n154 ) : ( n156 ) ;
assign n158 =  ( n153 ) ? ( 9'd0 ) : ( n157 ) ;
assign n159 =  ( n20 ) ? ( LB2D_shift_x ) : ( n158 ) ;
assign n160 =  ( n11 ) ? ( LB2D_shift_x ) : ( n159 ) ;
assign n161 =  ( n6 ) ? ( LB2D_shift_x ) : ( n160 ) ;
assign n162 =  ( LB2D_shift_y ) < ( 10'd640 )  ;
assign n163 =  ( LB2D_shift_x ) < ( 9'd488 )  ;
assign n164 =  ( LB2D_shift_y ) + ( 10'd1 )  ;
assign n165 =  ( n163 ) ? ( LB2D_shift_y ) : ( n164 ) ;
assign n166 =  ( n162 ) ? ( n165 ) : ( 10'd640 ) ;
assign n167 =  ( n39 ) ? ( LB2D_shift_y ) : ( LB2D_shift_y ) ;
assign n168 =  ( n34 ) ? ( LB2D_shift_y ) : ( n167 ) ;
assign n169 =  ( n29 ) ? ( n166 ) : ( n168 ) ;
assign n170 =  ( n20 ) ? ( LB2D_shift_y ) : ( n169 ) ;
assign n171 =  ( n11 ) ? ( LB2D_shift_y ) : ( n170 ) ;
assign n172 =  ( n6 ) ? ( LB2D_shift_y ) : ( n171 ) ;
assign n173 =  ( stencil_stream_full ) == ( 1'd1 )  ;
assign n174 =  ( n173 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_0 ) ;
assign n175 = gb_fun(n174) ;
assign n176 =  ( n39 ) ? ( arg_0_TDATA ) : ( arg_0_TDATA ) ;
assign n177 =  ( n34 ) ? ( arg_0_TDATA ) : ( n176 ) ;
assign n178 =  ( n29 ) ? ( arg_0_TDATA ) : ( n177 ) ;
assign n179 =  ( n20 ) ? ( n175 ) : ( n178 ) ;
assign n180 =  ( n11 ) ? ( arg_0_TDATA ) : ( n179 ) ;
assign n181 =  ( n6 ) ? ( arg_0_TDATA ) : ( n180 ) ;
assign n182 =  ( gb_pp_it_8 ) == ( 1'd1 )  ;
assign n183 =  ( n182 ) & ( n17 )  ;
assign n184 =  ( n183 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n185 =  ( n39 ) ? ( arg_0_TVALID ) : ( arg_0_TVALID ) ;
assign n186 =  ( n34 ) ? ( arg_0_TVALID ) : ( n185 ) ;
assign n187 =  ( n29 ) ? ( arg_0_TVALID ) : ( n186 ) ;
assign n188 =  ( n20 ) ? ( n184 ) : ( n187 ) ;
assign n189 =  ( n11 ) ? ( 1'd0 ) : ( n188 ) ;
assign n190 =  ( n6 ) ? ( arg_0_TVALID ) : ( n189 ) ;
assign n191 =  ( n39 ) ? ( 1'd1 ) : ( arg_1_TREADY ) ;
assign n192 =  ( n38 ) ? ( 1'd1 ) : ( n191 ) ;
assign n193 =  ( n34 ) ? ( arg_1_TREADY ) : ( n192 ) ;
assign n194 =  ( n29 ) ? ( arg_1_TREADY ) : ( n193 ) ;
assign n195 =  ( n20 ) ? ( arg_1_TREADY ) : ( n194 ) ;
assign n196 =  ( n11 ) ? ( arg_1_TREADY ) : ( n195 ) ;
assign n197 =  ( n6 ) ? ( 1'd1 ) : ( n196 ) ;
assign n198 =  ( gb_p_cnt ) == ( 19'd307200 )  ;
assign n199 =  ( n198 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n200 =  ( n39 ) ? ( gb_exit_it_1 ) : ( gb_exit_it_1 ) ;
assign n201 =  ( n34 ) ? ( gb_exit_it_1 ) : ( n200 ) ;
assign n202 =  ( n29 ) ? ( gb_exit_it_1 ) : ( n201 ) ;
assign n203 =  ( n20 ) ? ( n199 ) : ( n202 ) ;
assign n204 =  ( n11 ) ? ( gb_exit_it_1 ) : ( n203 ) ;
assign n205 =  ( n6 ) ? ( gb_exit_it_1 ) : ( n204 ) ;
assign n206 =  ( n39 ) ? ( gb_exit_it_2 ) : ( gb_exit_it_2 ) ;
assign n207 =  ( n34 ) ? ( gb_exit_it_2 ) : ( n206 ) ;
assign n208 =  ( n29 ) ? ( gb_exit_it_2 ) : ( n207 ) ;
assign n209 =  ( n20 ) ? ( gb_exit_it_1 ) : ( n208 ) ;
assign n210 =  ( n11 ) ? ( gb_exit_it_2 ) : ( n209 ) ;
assign n211 =  ( n6 ) ? ( gb_exit_it_2 ) : ( n210 ) ;
assign n212 =  ( n39 ) ? ( gb_exit_it_3 ) : ( gb_exit_it_3 ) ;
assign n213 =  ( n34 ) ? ( gb_exit_it_3 ) : ( n212 ) ;
assign n214 =  ( n29 ) ? ( gb_exit_it_3 ) : ( n213 ) ;
assign n215 =  ( n20 ) ? ( gb_exit_it_2 ) : ( n214 ) ;
assign n216 =  ( n11 ) ? ( gb_exit_it_3 ) : ( n215 ) ;
assign n217 =  ( n6 ) ? ( gb_exit_it_3 ) : ( n216 ) ;
assign n218 =  ( n39 ) ? ( gb_exit_it_4 ) : ( gb_exit_it_4 ) ;
assign n219 =  ( n34 ) ? ( gb_exit_it_4 ) : ( n218 ) ;
assign n220 =  ( n29 ) ? ( gb_exit_it_4 ) : ( n219 ) ;
assign n221 =  ( n20 ) ? ( gb_exit_it_3 ) : ( n220 ) ;
assign n222 =  ( n11 ) ? ( gb_exit_it_4 ) : ( n221 ) ;
assign n223 =  ( n6 ) ? ( gb_exit_it_4 ) : ( n222 ) ;
assign n224 =  ( n39 ) ? ( gb_exit_it_5 ) : ( gb_exit_it_5 ) ;
assign n225 =  ( n34 ) ? ( gb_exit_it_5 ) : ( n224 ) ;
assign n226 =  ( n29 ) ? ( gb_exit_it_5 ) : ( n225 ) ;
assign n227 =  ( n20 ) ? ( gb_exit_it_4 ) : ( n226 ) ;
assign n228 =  ( n11 ) ? ( gb_exit_it_5 ) : ( n227 ) ;
assign n229 =  ( n6 ) ? ( gb_exit_it_5 ) : ( n228 ) ;
assign n230 =  ( n39 ) ? ( gb_exit_it_6 ) : ( gb_exit_it_6 ) ;
assign n231 =  ( n34 ) ? ( gb_exit_it_6 ) : ( n230 ) ;
assign n232 =  ( n29 ) ? ( gb_exit_it_6 ) : ( n231 ) ;
assign n233 =  ( n20 ) ? ( gb_exit_it_5 ) : ( n232 ) ;
assign n234 =  ( n11 ) ? ( gb_exit_it_6 ) : ( n233 ) ;
assign n235 =  ( n6 ) ? ( gb_exit_it_6 ) : ( n234 ) ;
assign n236 =  ( n39 ) ? ( gb_exit_it_7 ) : ( gb_exit_it_7 ) ;
assign n237 =  ( n34 ) ? ( gb_exit_it_7 ) : ( n236 ) ;
assign n238 =  ( n29 ) ? ( gb_exit_it_7 ) : ( n237 ) ;
assign n239 =  ( n20 ) ? ( gb_exit_it_6 ) : ( n238 ) ;
assign n240 =  ( n11 ) ? ( gb_exit_it_7 ) : ( n239 ) ;
assign n241 =  ( n6 ) ? ( gb_exit_it_7 ) : ( n240 ) ;
assign n242 =  ( n39 ) ? ( gb_exit_it_8 ) : ( gb_exit_it_8 ) ;
assign n243 =  ( n34 ) ? ( gb_exit_it_8 ) : ( n242 ) ;
assign n244 =  ( n29 ) ? ( gb_exit_it_8 ) : ( n243 ) ;
assign n245 =  ( n20 ) ? ( gb_exit_it_7 ) : ( n244 ) ;
assign n246 =  ( n11 ) ? ( gb_exit_it_8 ) : ( n245 ) ;
assign n247 =  ( n6 ) ? ( gb_exit_it_8 ) : ( n246 ) ;
assign n248 =  ( gb_p_cnt ) < ( 19'd307200 )  ;
assign n249 =  ( gb_p_cnt ) + ( 19'd1 )  ;
assign n250 =  ( n248 ) ? ( n249 ) : ( 19'd307200 ) ;
assign n251 =  ( n39 ) ? ( gb_p_cnt ) : ( gb_p_cnt ) ;
assign n252 =  ( n34 ) ? ( gb_p_cnt ) : ( n251 ) ;
assign n253 =  ( n29 ) ? ( gb_p_cnt ) : ( n252 ) ;
assign n254 =  ( n20 ) ? ( n250 ) : ( n253 ) ;
assign n255 =  ( n11 ) ? ( gb_p_cnt ) : ( n254 ) ;
assign n256 =  ( n6 ) ? ( gb_p_cnt ) : ( n255 ) ;
assign n257 =  ( n39 ) ? ( gb_pp_it_1 ) : ( gb_pp_it_1 ) ;
assign n258 =  ( n34 ) ? ( gb_pp_it_1 ) : ( n257 ) ;
assign n259 =  ( n29 ) ? ( gb_pp_it_1 ) : ( n258 ) ;
assign n260 =  ( n20 ) ? ( 1'd1 ) : ( n259 ) ;
assign n261 =  ( n11 ) ? ( gb_pp_it_1 ) : ( n260 ) ;
assign n262 =  ( n6 ) ? ( gb_pp_it_1 ) : ( n261 ) ;
assign n263 =  ( n39 ) ? ( gb_pp_it_2 ) : ( gb_pp_it_2 ) ;
assign n264 =  ( n34 ) ? ( gb_pp_it_2 ) : ( n263 ) ;
assign n265 =  ( n29 ) ? ( gb_pp_it_2 ) : ( n264 ) ;
assign n266 =  ( n20 ) ? ( gb_pp_it_1 ) : ( n265 ) ;
assign n267 =  ( n11 ) ? ( gb_pp_it_2 ) : ( n266 ) ;
assign n268 =  ( n6 ) ? ( gb_pp_it_2 ) : ( n267 ) ;
assign n269 =  ( n39 ) ? ( gb_pp_it_3 ) : ( gb_pp_it_3 ) ;
assign n270 =  ( n34 ) ? ( gb_pp_it_3 ) : ( n269 ) ;
assign n271 =  ( n29 ) ? ( gb_pp_it_3 ) : ( n270 ) ;
assign n272 =  ( n20 ) ? ( gb_pp_it_2 ) : ( n271 ) ;
assign n273 =  ( n11 ) ? ( gb_pp_it_3 ) : ( n272 ) ;
assign n274 =  ( n6 ) ? ( gb_pp_it_3 ) : ( n273 ) ;
assign n275 =  ( n39 ) ? ( gb_pp_it_4 ) : ( gb_pp_it_4 ) ;
assign n276 =  ( n34 ) ? ( gb_pp_it_4 ) : ( n275 ) ;
assign n277 =  ( n29 ) ? ( gb_pp_it_4 ) : ( n276 ) ;
assign n278 =  ( n20 ) ? ( gb_pp_it_3 ) : ( n277 ) ;
assign n279 =  ( n11 ) ? ( gb_pp_it_4 ) : ( n278 ) ;
assign n280 =  ( n6 ) ? ( gb_pp_it_4 ) : ( n279 ) ;
assign n281 =  ( n39 ) ? ( gb_pp_it_5 ) : ( gb_pp_it_5 ) ;
assign n282 =  ( n34 ) ? ( gb_pp_it_5 ) : ( n281 ) ;
assign n283 =  ( n29 ) ? ( gb_pp_it_5 ) : ( n282 ) ;
assign n284 =  ( n20 ) ? ( gb_pp_it_4 ) : ( n283 ) ;
assign n285 =  ( n11 ) ? ( gb_pp_it_5 ) : ( n284 ) ;
assign n286 =  ( n6 ) ? ( gb_pp_it_5 ) : ( n285 ) ;
assign n287 =  ( n39 ) ? ( gb_pp_it_6 ) : ( gb_pp_it_6 ) ;
assign n288 =  ( n34 ) ? ( gb_pp_it_6 ) : ( n287 ) ;
assign n289 =  ( n29 ) ? ( gb_pp_it_6 ) : ( n288 ) ;
assign n290 =  ( n20 ) ? ( gb_pp_it_5 ) : ( n289 ) ;
assign n291 =  ( n11 ) ? ( gb_pp_it_6 ) : ( n290 ) ;
assign n292 =  ( n6 ) ? ( gb_pp_it_6 ) : ( n291 ) ;
assign n293 =  ( n39 ) ? ( gb_pp_it_7 ) : ( gb_pp_it_7 ) ;
assign n294 =  ( n34 ) ? ( gb_pp_it_7 ) : ( n293 ) ;
assign n295 =  ( n29 ) ? ( gb_pp_it_7 ) : ( n294 ) ;
assign n296 =  ( n20 ) ? ( gb_pp_it_6 ) : ( n295 ) ;
assign n297 =  ( n11 ) ? ( gb_pp_it_7 ) : ( n296 ) ;
assign n298 =  ( n6 ) ? ( gb_pp_it_7 ) : ( n297 ) ;
assign n299 =  ( n39 ) ? ( gb_pp_it_8 ) : ( gb_pp_it_8 ) ;
assign n300 =  ( n34 ) ? ( gb_pp_it_8 ) : ( n299 ) ;
assign n301 =  ( n29 ) ? ( gb_pp_it_8 ) : ( n300 ) ;
assign n302 =  ( n20 ) ? ( gb_pp_it_7 ) : ( n301 ) ;
assign n303 =  ( n11 ) ? ( gb_pp_it_8 ) : ( n302 ) ;
assign n304 =  ( n6 ) ? ( gb_pp_it_8 ) : ( n303 ) ;
assign n305 =  ( n39 ) ? ( gb_pp_it_9 ) : ( gb_pp_it_9 ) ;
assign n306 =  ( n34 ) ? ( gb_pp_it_9 ) : ( n305 ) ;
assign n307 =  ( n29 ) ? ( gb_pp_it_9 ) : ( n306 ) ;
assign n308 =  ( n20 ) ? ( gb_pp_it_8 ) : ( n307 ) ;
assign n309 =  ( n11 ) ? ( gb_pp_it_9 ) : ( n308 ) ;
assign n310 =  ( n6 ) ? ( gb_pp_it_9 ) : ( n309 ) ;
assign n311 =  ( n39 ) ? ( LB1D_uIn ) : ( in_stream_buff_0 ) ;
assign n312 =  ( n34 ) ? ( in_stream_buff_0 ) : ( n311 ) ;
assign n313 =  ( n29 ) ? ( in_stream_buff_0 ) : ( n312 ) ;
assign n314 =  ( n20 ) ? ( in_stream_buff_0 ) : ( n313 ) ;
assign n315 =  ( n11 ) ? ( in_stream_buff_0 ) : ( n314 ) ;
assign n316 =  ( n6 ) ? ( LB1D_uIn ) : ( n315 ) ;
assign n317 =  ( n39 ) ? ( in_stream_buff_0 ) : ( in_stream_buff_1 ) ;
assign n318 =  ( n34 ) ? ( in_stream_buff_1 ) : ( n317 ) ;
assign n319 =  ( n29 ) ? ( in_stream_buff_1 ) : ( n318 ) ;
assign n320 =  ( n20 ) ? ( in_stream_buff_1 ) : ( n319 ) ;
assign n321 =  ( n11 ) ? ( in_stream_buff_1 ) : ( n320 ) ;
assign n322 =  ( n6 ) ? ( in_stream_buff_0 ) : ( n321 ) ;
assign n323 =  ( in_stream_full ) == ( 1'd1 )  ;
assign n324 =  ( n323 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n325 =  ( n39 ) ? ( 1'd0 ) : ( in_stream_empty ) ;
assign n326 =  ( n34 ) ? ( n324 ) : ( n325 ) ;
assign n327 =  ( n29 ) ? ( in_stream_empty ) : ( n326 ) ;
assign n328 =  ( n20 ) ? ( in_stream_empty ) : ( n327 ) ;
assign n329 =  ( n11 ) ? ( in_stream_empty ) : ( n328 ) ;
assign n330 =  ( n6 ) ? ( 1'd0 ) : ( n329 ) ;
assign n331 =  ( in_stream_empty ) == ( 1'd1 )  ;
assign n332 =  ( n331 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n333 =  ( n39 ) ? ( n332 ) : ( in_stream_full ) ;
assign n334 =  ( n34 ) ? ( 1'd0 ) : ( n333 ) ;
assign n335 =  ( n29 ) ? ( in_stream_full ) : ( n334 ) ;
assign n336 =  ( n20 ) ? ( in_stream_full ) : ( n335 ) ;
assign n337 =  ( n11 ) ? ( in_stream_full ) : ( n336 ) ;
assign n338 =  ( n6 ) ? ( n332 ) : ( n337 ) ;
assign n339 =  ( n323 ) ? ( in_stream_buff_1 ) : ( in_stream_buff_0 ) ;
assign n340 =  ( LB2D_proc_w ) == ( 64'd0 )  ;
assign n341 =  ( LB2D_proc_x ) - ( 9'd1 )  ;
assign n342 =  (  LB2D_proc_7 [ n341 ] )  ;
assign n343 =  ( LB2D_proc_w ) == ( 64'd1 )  ;
assign n344 =  (  LB2D_proc_0 [ n341 ] )  ;
assign n345 =  ( LB2D_proc_w ) == ( 64'd2 )  ;
assign n346 =  (  LB2D_proc_1 [ n341 ] )  ;
assign n347 =  ( LB2D_proc_w ) == ( 64'd3 )  ;
assign n348 =  (  LB2D_proc_2 [ n341 ] )  ;
assign n349 =  ( LB2D_proc_w ) == ( 64'd4 )  ;
assign n350 =  (  LB2D_proc_3 [ n341 ] )  ;
assign n351 =  ( LB2D_proc_w ) == ( 64'd5 )  ;
assign n352 =  (  LB2D_proc_4 [ n341 ] )  ;
assign n353 =  ( LB2D_proc_w ) == ( 64'd6 )  ;
assign n354 =  (  LB2D_proc_5 [ n341 ] )  ;
assign n355 =  (  LB2D_proc_6 [ n341 ] )  ;
assign n356 =  ( n353 ) ? ( n354 ) : ( n355 ) ;
assign n357 =  ( n351 ) ? ( n352 ) : ( n356 ) ;
assign n358 =  ( n349 ) ? ( n350 ) : ( n357 ) ;
assign n359 =  ( n347 ) ? ( n348 ) : ( n358 ) ;
assign n360 =  ( n345 ) ? ( n346 ) : ( n359 ) ;
assign n361 =  ( n343 ) ? ( n344 ) : ( n360 ) ;
assign n362 =  ( n340 ) ? ( n342 ) : ( n361 ) ;
assign n363 =  ( n353 ) ? ( n352 ) : ( n354 ) ;
assign n364 =  ( n351 ) ? ( n350 ) : ( n363 ) ;
assign n365 =  ( n349 ) ? ( n348 ) : ( n364 ) ;
assign n366 =  ( n347 ) ? ( n346 ) : ( n365 ) ;
assign n367 =  ( n345 ) ? ( n344 ) : ( n366 ) ;
assign n368 =  ( n343 ) ? ( n342 ) : ( n367 ) ;
assign n369 =  ( n340 ) ? ( n355 ) : ( n368 ) ;
assign n370 =  ( n353 ) ? ( n350 ) : ( n352 ) ;
assign n371 =  ( n351 ) ? ( n348 ) : ( n370 ) ;
assign n372 =  ( n349 ) ? ( n346 ) : ( n371 ) ;
assign n373 =  ( n347 ) ? ( n344 ) : ( n372 ) ;
assign n374 =  ( n345 ) ? ( n342 ) : ( n373 ) ;
assign n375 =  ( n343 ) ? ( n355 ) : ( n374 ) ;
assign n376 =  ( n340 ) ? ( n354 ) : ( n375 ) ;
assign n377 =  ( n353 ) ? ( n348 ) : ( n350 ) ;
assign n378 =  ( n351 ) ? ( n346 ) : ( n377 ) ;
assign n379 =  ( n349 ) ? ( n344 ) : ( n378 ) ;
assign n380 =  ( n347 ) ? ( n342 ) : ( n379 ) ;
assign n381 =  ( n345 ) ? ( n355 ) : ( n380 ) ;
assign n382 =  ( n343 ) ? ( n354 ) : ( n381 ) ;
assign n383 =  ( n340 ) ? ( n352 ) : ( n382 ) ;
assign n384 =  ( n353 ) ? ( n346 ) : ( n348 ) ;
assign n385 =  ( n351 ) ? ( n344 ) : ( n384 ) ;
assign n386 =  ( n349 ) ? ( n342 ) : ( n385 ) ;
assign n387 =  ( n347 ) ? ( n355 ) : ( n386 ) ;
assign n388 =  ( n345 ) ? ( n354 ) : ( n387 ) ;
assign n389 =  ( n343 ) ? ( n352 ) : ( n388 ) ;
assign n390 =  ( n340 ) ? ( n350 ) : ( n389 ) ;
assign n391 =  ( n353 ) ? ( n344 ) : ( n346 ) ;
assign n392 =  ( n351 ) ? ( n342 ) : ( n391 ) ;
assign n393 =  ( n349 ) ? ( n355 ) : ( n392 ) ;
assign n394 =  ( n347 ) ? ( n354 ) : ( n393 ) ;
assign n395 =  ( n345 ) ? ( n352 ) : ( n394 ) ;
assign n396 =  ( n343 ) ? ( n350 ) : ( n395 ) ;
assign n397 =  ( n340 ) ? ( n348 ) : ( n396 ) ;
assign n398 =  ( n353 ) ? ( n342 ) : ( n344 ) ;
assign n399 =  ( n351 ) ? ( n355 ) : ( n398 ) ;
assign n400 =  ( n349 ) ? ( n354 ) : ( n399 ) ;
assign n401 =  ( n347 ) ? ( n352 ) : ( n400 ) ;
assign n402 =  ( n345 ) ? ( n350 ) : ( n401 ) ;
assign n403 =  ( n343 ) ? ( n348 ) : ( n402 ) ;
assign n404 =  ( n340 ) ? ( n346 ) : ( n403 ) ;
assign n405 =  ( n353 ) ? ( n355 ) : ( n342 ) ;
assign n406 =  ( n351 ) ? ( n354 ) : ( n405 ) ;
assign n407 =  ( n349 ) ? ( n352 ) : ( n406 ) ;
assign n408 =  ( n347 ) ? ( n350 ) : ( n407 ) ;
assign n409 =  ( n345 ) ? ( n348 ) : ( n408 ) ;
assign n410 =  ( n343 ) ? ( n346 ) : ( n409 ) ;
assign n411 =  ( n340 ) ? ( n344 ) : ( n410 ) ;
assign n412 =  { ( n404 ) , ( n411 ) }  ;
assign n413 =  { ( n397 ) , ( n412 ) }  ;
assign n414 =  { ( n390 ) , ( n413 ) }  ;
assign n415 =  { ( n383 ) , ( n414 ) }  ;
assign n416 =  { ( n376 ) , ( n415 ) }  ;
assign n417 =  { ( n369 ) , ( n416 ) }  ;
assign n418 =  { ( n362 ) , ( n417 ) }  ;
assign n419 =  { ( n339 ) , ( n418 ) }  ;
assign n420 =  ( n32 ) ? ( slice_stream_buff_0 ) : ( n419 ) ;
assign n421 =  ( n39 ) ? ( slice_stream_buff_0 ) : ( slice_stream_buff_0 ) ;
assign n422 =  ( n34 ) ? ( n420 ) : ( n421 ) ;
assign n423 =  ( n29 ) ? ( slice_stream_buff_0 ) : ( n422 ) ;
assign n424 =  ( n20 ) ? ( slice_stream_buff_0 ) : ( n423 ) ;
assign n425 =  ( n11 ) ? ( slice_stream_buff_0 ) : ( n424 ) ;
assign n426 =  ( n6 ) ? ( slice_stream_buff_0 ) : ( n425 ) ;
assign n427 =  ( n32 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n428 =  ( n39 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_1 ) ;
assign n429 =  ( n34 ) ? ( n427 ) : ( n428 ) ;
assign n430 =  ( n29 ) ? ( slice_stream_buff_1 ) : ( n429 ) ;
assign n431 =  ( n20 ) ? ( slice_stream_buff_1 ) : ( n430 ) ;
assign n432 =  ( n11 ) ? ( slice_stream_buff_1 ) : ( n431 ) ;
assign n433 =  ( n6 ) ? ( slice_stream_buff_1 ) : ( n432 ) ;
assign n434 =  ( n142 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n435 =  ( n32 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n436 =  ( n39 ) ? ( slice_stream_empty ) : ( slice_stream_empty ) ;
assign n437 =  ( n34 ) ? ( n435 ) : ( n436 ) ;
assign n438 =  ( n29 ) ? ( n434 ) : ( n437 ) ;
assign n439 =  ( n20 ) ? ( slice_stream_empty ) : ( n438 ) ;
assign n440 =  ( n11 ) ? ( slice_stream_empty ) : ( n439 ) ;
assign n441 =  ( n6 ) ? ( slice_stream_empty ) : ( n440 ) ;
assign n442 =  ( slice_stream_empty ) == ( 1'd1 )  ;
assign n443 =  ( n442 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n444 =  ( n32 ) ? ( 1'd0 ) : ( n443 ) ;
assign n445 =  ( n39 ) ? ( slice_stream_full ) : ( slice_stream_full ) ;
assign n446 =  ( n34 ) ? ( n444 ) : ( n445 ) ;
assign n447 =  ( n29 ) ? ( 1'd0 ) : ( n446 ) ;
assign n448 =  ( n20 ) ? ( slice_stream_full ) : ( n447 ) ;
assign n449 =  ( n11 ) ? ( slice_stream_full ) : ( n448 ) ;
assign n450 =  ( n6 ) ? ( slice_stream_full ) : ( n449 ) ;
assign n451 =  ( LB2D_shift_x ) >= ( 9'd8 )  ;
assign n452 =  ( LB2D_shift_x ) == ( 9'd0 )  ;
assign n453 =  ( n451 ) | ( n452 )  ;
assign n454 = n143[71:64] ;
assign n455 = LB2D_shift_7[71:64] ;
assign n456 = LB2D_shift_6[71:64] ;
assign n457 = LB2D_shift_5[71:64] ;
assign n458 = LB2D_shift_4[71:64] ;
assign n459 = LB2D_shift_3[71:64] ;
assign n460 = LB2D_shift_2[71:64] ;
assign n461 = LB2D_shift_1[71:64] ;
assign n462 = LB2D_shift_0[71:64] ;
assign n463 =  { ( n461 ) , ( n462 ) }  ;
assign n464 =  { ( n460 ) , ( n463 ) }  ;
assign n465 =  { ( n459 ) , ( n464 ) }  ;
assign n466 =  { ( n458 ) , ( n465 ) }  ;
assign n467 =  { ( n457 ) , ( n466 ) }  ;
assign n468 =  { ( n456 ) , ( n467 ) }  ;
assign n469 =  { ( n455 ) , ( n468 ) }  ;
assign n470 =  { ( n454 ) , ( n469 ) }  ;
assign n471 = n143[63:56] ;
assign n472 = LB2D_shift_7[63:56] ;
assign n473 = LB2D_shift_6[63:56] ;
assign n474 = LB2D_shift_5[63:56] ;
assign n475 = LB2D_shift_4[63:56] ;
assign n476 = LB2D_shift_3[63:56] ;
assign n477 = LB2D_shift_2[63:56] ;
assign n478 = LB2D_shift_1[63:56] ;
assign n479 = LB2D_shift_0[63:56] ;
assign n480 =  { ( n478 ) , ( n479 ) }  ;
assign n481 =  { ( n477 ) , ( n480 ) }  ;
assign n482 =  { ( n476 ) , ( n481 ) }  ;
assign n483 =  { ( n475 ) , ( n482 ) }  ;
assign n484 =  { ( n474 ) , ( n483 ) }  ;
assign n485 =  { ( n473 ) , ( n484 ) }  ;
assign n486 =  { ( n472 ) , ( n485 ) }  ;
assign n487 =  { ( n471 ) , ( n486 ) }  ;
assign n488 = n143[55:48] ;
assign n489 = LB2D_shift_7[55:48] ;
assign n490 = LB2D_shift_6[55:48] ;
assign n491 = LB2D_shift_5[55:48] ;
assign n492 = LB2D_shift_4[55:48] ;
assign n493 = LB2D_shift_3[55:48] ;
assign n494 = LB2D_shift_2[55:48] ;
assign n495 = LB2D_shift_1[55:48] ;
assign n496 = LB2D_shift_0[55:48] ;
assign n497 =  { ( n495 ) , ( n496 ) }  ;
assign n498 =  { ( n494 ) , ( n497 ) }  ;
assign n499 =  { ( n493 ) , ( n498 ) }  ;
assign n500 =  { ( n492 ) , ( n499 ) }  ;
assign n501 =  { ( n491 ) , ( n500 ) }  ;
assign n502 =  { ( n490 ) , ( n501 ) }  ;
assign n503 =  { ( n489 ) , ( n502 ) }  ;
assign n504 =  { ( n488 ) , ( n503 ) }  ;
assign n505 = n143[47:40] ;
assign n506 = LB2D_shift_7[47:40] ;
assign n507 = LB2D_shift_6[47:40] ;
assign n508 = LB2D_shift_5[47:40] ;
assign n509 = LB2D_shift_4[47:40] ;
assign n510 = LB2D_shift_3[47:40] ;
assign n511 = LB2D_shift_2[47:40] ;
assign n512 = LB2D_shift_1[47:40] ;
assign n513 = LB2D_shift_0[47:40] ;
assign n514 =  { ( n512 ) , ( n513 ) }  ;
assign n515 =  { ( n511 ) , ( n514 ) }  ;
assign n516 =  { ( n510 ) , ( n515 ) }  ;
assign n517 =  { ( n509 ) , ( n516 ) }  ;
assign n518 =  { ( n508 ) , ( n517 ) }  ;
assign n519 =  { ( n507 ) , ( n518 ) }  ;
assign n520 =  { ( n506 ) , ( n519 ) }  ;
assign n521 =  { ( n505 ) , ( n520 ) }  ;
assign n522 = n143[39:32] ;
assign n523 = LB2D_shift_7[39:32] ;
assign n524 = LB2D_shift_6[39:32] ;
assign n525 = LB2D_shift_5[39:32] ;
assign n526 = LB2D_shift_4[39:32] ;
assign n527 = LB2D_shift_3[39:32] ;
assign n528 = LB2D_shift_2[39:32] ;
assign n529 = LB2D_shift_1[39:32] ;
assign n530 = LB2D_shift_0[39:32] ;
assign n531 =  { ( n529 ) , ( n530 ) }  ;
assign n532 =  { ( n528 ) , ( n531 ) }  ;
assign n533 =  { ( n527 ) , ( n532 ) }  ;
assign n534 =  { ( n526 ) , ( n533 ) }  ;
assign n535 =  { ( n525 ) , ( n534 ) }  ;
assign n536 =  { ( n524 ) , ( n535 ) }  ;
assign n537 =  { ( n523 ) , ( n536 ) }  ;
assign n538 =  { ( n522 ) , ( n537 ) }  ;
assign n539 = n143[31:24] ;
assign n540 = LB2D_shift_7[31:24] ;
assign n541 = LB2D_shift_6[31:24] ;
assign n542 = LB2D_shift_5[31:24] ;
assign n543 = LB2D_shift_4[31:24] ;
assign n544 = LB2D_shift_3[31:24] ;
assign n545 = LB2D_shift_2[31:24] ;
assign n546 = LB2D_shift_1[31:24] ;
assign n547 = LB2D_shift_0[31:24] ;
assign n548 =  { ( n546 ) , ( n547 ) }  ;
assign n549 =  { ( n545 ) , ( n548 ) }  ;
assign n550 =  { ( n544 ) , ( n549 ) }  ;
assign n551 =  { ( n543 ) , ( n550 ) }  ;
assign n552 =  { ( n542 ) , ( n551 ) }  ;
assign n553 =  { ( n541 ) , ( n552 ) }  ;
assign n554 =  { ( n540 ) , ( n553 ) }  ;
assign n555 =  { ( n539 ) , ( n554 ) }  ;
assign n556 = n143[23:16] ;
assign n557 = LB2D_shift_7[23:16] ;
assign n558 = LB2D_shift_6[23:16] ;
assign n559 = LB2D_shift_5[23:16] ;
assign n560 = LB2D_shift_4[23:16] ;
assign n561 = LB2D_shift_3[23:16] ;
assign n562 = LB2D_shift_2[23:16] ;
assign n563 = LB2D_shift_1[23:16] ;
assign n564 = LB2D_shift_0[23:16] ;
assign n565 =  { ( n563 ) , ( n564 ) }  ;
assign n566 =  { ( n562 ) , ( n565 ) }  ;
assign n567 =  { ( n561 ) , ( n566 ) }  ;
assign n568 =  { ( n560 ) , ( n567 ) }  ;
assign n569 =  { ( n559 ) , ( n568 ) }  ;
assign n570 =  { ( n558 ) , ( n569 ) }  ;
assign n571 =  { ( n557 ) , ( n570 ) }  ;
assign n572 =  { ( n556 ) , ( n571 ) }  ;
assign n573 = n143[15:8] ;
assign n574 = LB2D_shift_7[15:8] ;
assign n575 = LB2D_shift_6[15:8] ;
assign n576 = LB2D_shift_5[15:8] ;
assign n577 = LB2D_shift_4[15:8] ;
assign n578 = LB2D_shift_3[15:8] ;
assign n579 = LB2D_shift_2[15:8] ;
assign n580 = LB2D_shift_1[15:8] ;
assign n581 = LB2D_shift_0[15:8] ;
assign n582 =  { ( n580 ) , ( n581 ) }  ;
assign n583 =  { ( n579 ) , ( n582 ) }  ;
assign n584 =  { ( n578 ) , ( n583 ) }  ;
assign n585 =  { ( n577 ) , ( n584 ) }  ;
assign n586 =  { ( n576 ) , ( n585 ) }  ;
assign n587 =  { ( n575 ) , ( n586 ) }  ;
assign n588 =  { ( n574 ) , ( n587 ) }  ;
assign n589 =  { ( n573 ) , ( n588 ) }  ;
assign n590 = n143[7:0] ;
assign n591 = LB2D_shift_7[7:0] ;
assign n592 = LB2D_shift_6[7:0] ;
assign n593 = LB2D_shift_5[7:0] ;
assign n594 = LB2D_shift_4[7:0] ;
assign n595 = LB2D_shift_3[7:0] ;
assign n596 = LB2D_shift_2[7:0] ;
assign n597 = LB2D_shift_1[7:0] ;
assign n598 = LB2D_shift_0[7:0] ;
assign n599 =  { ( n597 ) , ( n598 ) }  ;
assign n600 =  { ( n596 ) , ( n599 ) }  ;
assign n601 =  { ( n595 ) , ( n600 ) }  ;
assign n602 =  { ( n594 ) , ( n601 ) }  ;
assign n603 =  { ( n593 ) , ( n602 ) }  ;
assign n604 =  { ( n592 ) , ( n603 ) }  ;
assign n605 =  { ( n591 ) , ( n604 ) }  ;
assign n606 =  { ( n590 ) , ( n605 ) }  ;
assign n607 =  { ( n589 ) , ( n606 ) }  ;
assign n608 =  { ( n572 ) , ( n607 ) }  ;
assign n609 =  { ( n555 ) , ( n608 ) }  ;
assign n610 =  { ( n538 ) , ( n609 ) }  ;
assign n611 =  { ( n521 ) , ( n610 ) }  ;
assign n612 =  { ( n504 ) , ( n611 ) }  ;
assign n613 =  { ( n487 ) , ( n612 ) }  ;
assign n614 =  { ( n470 ) , ( n613 ) }  ;
assign n615 =  ( n453 ) ? ( n614 ) : ( stencil_stream_buff_0 ) ;
assign n616 =  ( n39 ) ? ( stencil_stream_buff_0 ) : ( stencil_stream_buff_0 ) ;
assign n617 =  ( n34 ) ? ( stencil_stream_buff_0 ) : ( n616 ) ;
assign n618 =  ( n29 ) ? ( n615 ) : ( n617 ) ;
assign n619 =  ( n20 ) ? ( stencil_stream_buff_0 ) : ( n618 ) ;
assign n620 =  ( n11 ) ? ( stencil_stream_buff_0 ) : ( n619 ) ;
assign n621 =  ( n6 ) ? ( stencil_stream_buff_0 ) : ( n620 ) ;
assign n622 =  ( n39 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_1 ) ;
assign n623 =  ( n34 ) ? ( stencil_stream_buff_1 ) : ( n622 ) ;
assign n624 =  ( n29 ) ? ( stencil_stream_buff_0 ) : ( n623 ) ;
assign n625 =  ( n20 ) ? ( stencil_stream_buff_1 ) : ( n624 ) ;
assign n626 =  ( n11 ) ? ( stencil_stream_buff_1 ) : ( n625 ) ;
assign n627 =  ( n6 ) ? ( stencil_stream_buff_1 ) : ( n626 ) ;
assign n628 =  ( n173 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n629 = ~ ( n453 ) ;
assign n630 =  ( n629 ) ? ( stencil_stream_empty ) : ( 1'd0 ) ;
assign n631 =  ( n39 ) ? ( stencil_stream_empty ) : ( stencil_stream_empty ) ;
assign n632 =  ( n34 ) ? ( stencil_stream_empty ) : ( n631 ) ;
assign n633 =  ( n29 ) ? ( n630 ) : ( n632 ) ;
assign n634 =  ( n20 ) ? ( n628 ) : ( n633 ) ;
assign n635 =  ( n11 ) ? ( stencil_stream_empty ) : ( n634 ) ;
assign n636 =  ( n6 ) ? ( stencil_stream_empty ) : ( n635 ) ;
assign n637 =  ( n16 ) ? ( 1'd0 ) : ( 1'd0 ) ;
assign n638 =  ( stencil_stream_empty ) == ( 1'd1 )  ;
assign n639 =  ( n638 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n640 =  ( n629 ) ? ( stencil_stream_full ) : ( n639 ) ;
assign n641 =  ( n39 ) ? ( stencil_stream_full ) : ( stencil_stream_full ) ;
assign n642 =  ( n34 ) ? ( stencil_stream_full ) : ( n641 ) ;
assign n643 =  ( n29 ) ? ( n640 ) : ( n642 ) ;
assign n644 =  ( n20 ) ? ( n637 ) : ( n643 ) ;
assign n645 =  ( n11 ) ? ( stencil_stream_full ) : ( n644 ) ;
assign n646 =  ( n6 ) ? ( stencil_stream_full ) : ( n645 ) ;
assign n647 = ~ ( n6 ) ;
assign n648 = ~ ( n11 ) ;
assign n649 =  ( n647 ) & ( n648 )  ;
assign n650 = ~ ( n20 ) ;
assign n651 =  ( n649 ) & ( n650 )  ;
assign n652 = ~ ( n29 ) ;
assign n653 =  ( n651 ) & ( n652 )  ;
assign n654 = ~ ( n34 ) ;
assign n655 =  ( n653 ) & ( n654 )  ;
assign n656 = ~ ( n39 ) ;
assign n657 =  ( n655 ) & ( n656 )  ;
assign n658 =  ( n655 ) & ( n39 )  ;
assign n659 =  ( n653 ) & ( n34 )  ;
assign n660 = ~ ( n340 ) ;
assign n661 =  ( n659 ) & ( n660 )  ;
assign n662 =  ( n659 ) & ( n340 )  ;
assign n663 =  ( n651 ) & ( n29 )  ;
assign n664 =  ( n649 ) & ( n20 )  ;
assign n665 =  ( n647 ) & ( n11 )  ;
assign LB2D_proc_0_addr0 = n662 ? (n341) : (0);
assign LB2D_proc_0_data0 = n662 ? (n339) : (LB2D_proc_0[0]);
assign n666 = ~ ( n343 ) ;
assign n667 =  ( n659 ) & ( n666 )  ;
assign n668 =  ( n659 ) & ( n343 )  ;
assign LB2D_proc_1_addr0 = n668 ? (n341) : (0);
assign LB2D_proc_1_data0 = n668 ? (n339) : (LB2D_proc_1[0]);
assign n669 = ~ ( n345 ) ;
assign n670 =  ( n659 ) & ( n669 )  ;
assign n671 =  ( n659 ) & ( n345 )  ;
assign LB2D_proc_2_addr0 = n671 ? (n341) : (0);
assign LB2D_proc_2_data0 = n671 ? (n339) : (LB2D_proc_2[0]);
assign n672 = ~ ( n347 ) ;
assign n673 =  ( n659 ) & ( n672 )  ;
assign n674 =  ( n659 ) & ( n347 )  ;
assign LB2D_proc_3_addr0 = n674 ? (n341) : (0);
assign LB2D_proc_3_data0 = n674 ? (n339) : (LB2D_proc_3[0]);
assign n675 = ~ ( n349 ) ;
assign n676 =  ( n659 ) & ( n675 )  ;
assign n677 =  ( n659 ) & ( n349 )  ;
assign LB2D_proc_4_addr0 = n677 ? (n341) : (0);
assign LB2D_proc_4_data0 = n677 ? (n339) : (LB2D_proc_4[0]);
assign n678 = ~ ( n351 ) ;
assign n679 =  ( n659 ) & ( n678 )  ;
assign n680 =  ( n659 ) & ( n351 )  ;
assign LB2D_proc_5_addr0 = n680 ? (n341) : (0);
assign LB2D_proc_5_data0 = n680 ? (n339) : (LB2D_proc_5[0]);
assign n681 = ~ ( n353 ) ;
assign n682 =  ( n659 ) & ( n681 )  ;
assign n683 =  ( n659 ) & ( n353 )  ;
assign LB2D_proc_6_addr0 = n683 ? (n341) : (0);
assign LB2D_proc_6_data0 = n683 ? (n339) : (LB2D_proc_6[0]);
assign n684 = ~ ( n72 ) ;
assign n685 =  ( n659 ) & ( n684 )  ;
assign n686 =  ( n659 ) & ( n72 )  ;
assign LB2D_proc_7_addr0 = n686 ? (n341) : (0);
assign LB2D_proc_7_data0 = n686 ? (n339) : (LB2D_proc_7[0]);
/*
function [7:0] gb_fun ;
input [647:0] arg0;
    begin
//TODO: Add the specific function HERE.    end
endfunction
*/

always @(posedge clk) begin
   if(rst) begin
       LB1D_buff <= LB1D_buff;
       LB1D_in <= LB1D_in;
       LB1D_it_1 <= LB1D_it_1;
       LB1D_p_cnt <= LB1D_p_cnt;
       LB1D_uIn <= LB1D_uIn;
       LB2D_proc_w <= LB2D_proc_w;
       LB2D_proc_x <= LB2D_proc_x;
       LB2D_proc_y <= LB2D_proc_y;
       LB2D_shift_0 <= LB2D_shift_0;
       LB2D_shift_1 <= LB2D_shift_1;
       LB2D_shift_2 <= LB2D_shift_2;
       LB2D_shift_3 <= LB2D_shift_3;
       LB2D_shift_4 <= LB2D_shift_4;
       LB2D_shift_5 <= LB2D_shift_5;
       LB2D_shift_6 <= LB2D_shift_6;
       LB2D_shift_7 <= LB2D_shift_7;
       LB2D_shift_x <= LB2D_shift_x;
       LB2D_shift_y <= LB2D_shift_y;
       arg_0_TDATA <= arg_0_TDATA;
       arg_0_TVALID <= arg_0_TVALID;
       arg_1_TREADY <= arg_1_TREADY;
       gb_exit_it_1 <= gb_exit_it_1;
       gb_exit_it_2 <= gb_exit_it_2;
       gb_exit_it_3 <= gb_exit_it_3;
       gb_exit_it_4 <= gb_exit_it_4;
       gb_exit_it_5 <= gb_exit_it_5;
       gb_exit_it_6 <= gb_exit_it_6;
       gb_exit_it_7 <= gb_exit_it_7;
       gb_exit_it_8 <= gb_exit_it_8;
       gb_p_cnt <= gb_p_cnt;
       gb_pp_it_1 <= gb_pp_it_1;
       gb_pp_it_2 <= gb_pp_it_2;
       gb_pp_it_3 <= gb_pp_it_3;
       gb_pp_it_4 <= gb_pp_it_4;
       gb_pp_it_5 <= gb_pp_it_5;
       gb_pp_it_6 <= gb_pp_it_6;
       gb_pp_it_7 <= gb_pp_it_7;
       gb_pp_it_8 <= gb_pp_it_8;
       gb_pp_it_9 <= gb_pp_it_9;
       in_stream_buff_0 <= in_stream_buff_0;
       in_stream_buff_1 <= in_stream_buff_1;
       in_stream_empty <= in_stream_empty;
       in_stream_full <= in_stream_full;
       slice_stream_buff_0 <= slice_stream_buff_0;
       slice_stream_buff_1 <= slice_stream_buff_1;
       slice_stream_empty <= slice_stream_empty;
       slice_stream_full <= slice_stream_full;
       stencil_stream_buff_0 <= stencil_stream_buff_0;
       stencil_stream_buff_1 <= stencil_stream_buff_1;
       stencil_stream_empty <= stencil_stream_empty;
       stencil_stream_full <= stencil_stream_full;
   end
   else if(step) begin
       LB1D_buff <= n46;
       LB1D_in <= n53;
       LB1D_it_1 <= n56;
       LB1D_p_cnt <= n64;
       LB1D_uIn <= n70;
       LB2D_proc_w <= n81;
       LB2D_proc_x <= n89;
       LB2D_proc_y <= n99;
       LB2D_shift_0 <= n105;
       LB2D_shift_1 <= n111;
       LB2D_shift_2 <= n117;
       LB2D_shift_3 <= n123;
       LB2D_shift_4 <= n129;
       LB2D_shift_5 <= n135;
       LB2D_shift_6 <= n141;
       LB2D_shift_7 <= n149;
       LB2D_shift_x <= n161;
       LB2D_shift_y <= n172;
       arg_0_TDATA <= n181;
       arg_0_TVALID <= n190;
       arg_1_TREADY <= n197;
       gb_exit_it_1 <= n205;
       gb_exit_it_2 <= n211;
       gb_exit_it_3 <= n217;
       gb_exit_it_4 <= n223;
       gb_exit_it_5 <= n229;
       gb_exit_it_6 <= n235;
       gb_exit_it_7 <= n241;
       gb_exit_it_8 <= n247;
       gb_p_cnt <= n256;
       gb_pp_it_1 <= n262;
       gb_pp_it_2 <= n268;
       gb_pp_it_3 <= n274;
       gb_pp_it_4 <= n280;
       gb_pp_it_5 <= n286;
       gb_pp_it_6 <= n292;
       gb_pp_it_7 <= n298;
       gb_pp_it_8 <= n304;
       gb_pp_it_9 <= n310;
       in_stream_buff_0 <= n316;
       in_stream_buff_1 <= n322;
       in_stream_empty <= n330;
       in_stream_full <= n338;
       slice_stream_buff_0 <= n426;
       slice_stream_buff_1 <= n433;
       slice_stream_empty <= n441;
       slice_stream_full <= n450;
       stencil_stream_buff_0 <= n621;
       stencil_stream_buff_1 <= n627;
       stencil_stream_empty <= n636;
       stencil_stream_full <= n646;
       LB2D_proc_0 [ LB2D_proc_0_addr0 ] <= LB2D_proc_0_data0;
       LB2D_proc_1 [ LB2D_proc_1_addr0 ] <= LB2D_proc_1_data0;
       LB2D_proc_2 [ LB2D_proc_2_addr0 ] <= LB2D_proc_2_data0;
       LB2D_proc_3 [ LB2D_proc_3_addr0 ] <= LB2D_proc_3_data0;
       LB2D_proc_4 [ LB2D_proc_4_addr0 ] <= LB2D_proc_4_data0;
       LB2D_proc_5 [ LB2D_proc_5_addr0 ] <= LB2D_proc_5_data0;
       LB2D_proc_6 [ LB2D_proc_6_addr0 ] <= LB2D_proc_6_data0;
       LB2D_proc_7 [ LB2D_proc_7_addr0 ] <= LB2D_proc_7_data0;
   end
end
endmodule
