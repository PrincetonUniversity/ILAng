module ALU(
  input   clock,
  input   reset,
  input   io_dw,
  input  [3:0] io_fn,
  input  [31:0] io_in2,
  input  [31:0] io_in1,
  output [31:0] io_out,
  output [31:0] io_adder_out,
  output  io_cmp_out
);
  wire  T_15;
  wire [31:0] T_16;
  wire [31:0] in2_inv;
  wire [31:0] in1_xor_in2;
  wire [32:0] T_17;
  wire [31:0] T_18;
  wire [31:0] GEN_0;
  wire [32:0] T_20;
  wire [31:0] T_21;
  wire  T_22;
  wire  T_25;
  wire  T_27;
  wire  T_28;
  wire  T_29;
  wire  T_30;
  wire  T_31;
  wire  T_32;
  wire  T_35;
  wire  T_36;
  wire  T_37;
  wire  T_38;
  wire [4:0] shamt;
  wire  T_39;
  wire  T_40;
  wire  T_41;
  wire [15:0] T_46;
  wire [31:0] T_47;
  wire [15:0] T_48;
  wire [31:0] GEN_1;
  wire [31:0] T_49;
  wire [31:0] T_51;
  wire [31:0] T_52;
  wire [23:0] T_56;
  wire [31:0] GEN_2;
  wire [31:0] T_57;
  wire [23:0] T_58;
  wire [31:0] GEN_3;
  wire [31:0] T_59;
  wire [31:0] T_61;
  wire [31:0] T_62;
  wire [27:0] T_66;
  wire [31:0] GEN_4;
  wire [31:0] T_67;
  wire [27:0] T_68;
  wire [31:0] GEN_5;
  wire [31:0] T_69;
  wire [31:0] T_71;
  wire [31:0] T_72;
  wire [29:0] T_76;
  wire [31:0] GEN_6;
  wire [31:0] T_77;
  wire [29:0] T_78;
  wire [31:0] GEN_7;
  wire [31:0] T_79;
  wire [31:0] T_81;
  wire [31:0] T_82;
  wire [30:0] T_86;
  wire [31:0] GEN_8;
  wire [31:0] T_87;
  wire [30:0] T_88;
  wire [31:0] GEN_9;
  wire [31:0] T_89;
  wire [31:0] T_91;
  wire [31:0] T_92;
  wire [31:0] shin;
  wire  T_94;
  wire  T_95;
  wire [32:0] T_96;
  wire [32:0] T_97;
  wire [32:0] T_98;
  wire [31:0] shout_r;
  wire [15:0] T_103;
  wire [31:0] T_104;
  wire [15:0] T_105;
  wire [31:0] GEN_10;
  wire [31:0] T_106;
  wire [31:0] T_108;
  wire [31:0] T_109;
  wire [23:0] T_113;
  wire [31:0] GEN_11;
  wire [31:0] T_114;
  wire [23:0] T_115;
  wire [31:0] GEN_12;
  wire [31:0] T_116;
  wire [31:0] T_118;
  wire [31:0] T_119;
  wire [27:0] T_123;
  wire [31:0] GEN_13;
  wire [31:0] T_124;
  wire [27:0] T_125;
  wire [31:0] GEN_14;
  wire [31:0] T_126;
  wire [31:0] T_128;
  wire [31:0] T_129;
  wire [29:0] T_133;
  wire [31:0] GEN_15;
  wire [31:0] T_134;
  wire [29:0] T_135;
  wire [31:0] GEN_16;
  wire [31:0] T_136;
  wire [31:0] T_138;
  wire [31:0] T_139;
  wire [30:0] T_143;
  wire [31:0] GEN_17;
  wire [31:0] T_144;
  wire [30:0] T_145;
  wire [31:0] GEN_18;
  wire [31:0] T_146;
  wire [31:0] T_148;
  wire [31:0] shout_l;
  wire [31:0] T_153;
  wire  T_154;
  wire [31:0] T_156;
  wire [31:0] shout;
  wire  T_157;
  wire  T_158;
  wire  T_159;
  wire [31:0] T_161;
  wire  T_163;
  wire  T_164;
  wire [31:0] T_165;
  wire [31:0] T_167;
  wire [31:0] logic$;
  wire  T_168;
  wire  T_169;
  wire  T_170;
  wire  T_171;
  wire  T_172;
  wire  T_173;
  wire [31:0] GEN_19;
  wire [31:0] T_174;
  wire [31:0] shift_logic;
  wire  T_175;
  wire  T_176;
  wire  T_177;
  wire [31:0] out;
  assign io_out = out;
  assign io_adder_out = T_21;
  assign io_cmp_out = T_38;
  assign T_15 = io_fn[3];
  assign T_16 = ~ io_in2;
  assign in2_inv = T_15 ? T_16 : io_in2;
  assign in1_xor_in2 = io_in1 ^ in2_inv;
  assign T_17 = io_in1 + in2_inv;
  assign T_18 = T_17[31:0];
  assign GEN_0 = {{31'd0}, T_15};
  assign T_20 = T_18 + GEN_0;
  assign T_21 = T_20[31:0];
  assign T_22 = io_fn[0];
  assign T_25 = T_15 == 1'h0;
  assign T_27 = in1_xor_in2 == 32'h0;
  assign T_28 = io_in1[31];
  assign T_29 = io_in2[31];
  assign T_30 = T_28 == T_29;
  assign T_31 = io_adder_out[31];
  assign T_32 = io_fn[1];
  assign T_35 = T_32 ? T_29 : T_28;
  assign T_36 = T_30 ? T_31 : T_35;
  assign T_37 = T_25 ? T_27 : T_36;
  assign T_38 = T_22 ^ T_37;
  assign shamt = io_in2[4:0];
  assign T_39 = io_fn == 4'h5;
  assign T_40 = io_fn == 4'hb;
  assign T_41 = T_39 | T_40;
  assign T_46 = io_in1[31:16];
  assign T_47 = {{16'd0}, T_46};
  assign T_48 = io_in1[15:0];
  assign GEN_1 = {{16'd0}, T_48};
  assign T_49 = GEN_1 << 16;
  assign T_51 = T_49 & 32'hffff0000;
  assign T_52 = T_47 | T_51;
  assign T_56 = T_52[31:8];
  assign GEN_2 = {{8'd0}, T_56};
  assign T_57 = GEN_2 & 32'hff00ff;
  assign T_58 = T_52[23:0];
  assign GEN_3 = {{8'd0}, T_58};
  assign T_59 = GEN_3 << 8;
  assign T_61 = T_59 & 32'hff00ff00;
  assign T_62 = T_57 | T_61;
  assign T_66 = T_62[31:4];
  assign GEN_4 = {{4'd0}, T_66};
  assign T_67 = GEN_4 & 32'hf0f0f0f;
  assign T_68 = T_62[27:0];
  assign GEN_5 = {{4'd0}, T_68};
  assign T_69 = GEN_5 << 4;
  assign T_71 = T_69 & 32'hf0f0f0f0;
  assign T_72 = T_67 | T_71;
  assign T_76 = T_72[31:2];
  assign GEN_6 = {{2'd0}, T_76};
  assign T_77 = GEN_6 & 32'h33333333;
  assign T_78 = T_72[29:0];
  assign GEN_7 = {{2'd0}, T_78};
  assign T_79 = GEN_7 << 2;
  assign T_81 = T_79 & 32'hcccccccc;
  assign T_82 = T_77 | T_81;
  assign T_86 = T_82[31:1];
  assign GEN_8 = {{1'd0}, T_86};
  assign T_87 = GEN_8 & 32'h55555555;
  assign T_88 = T_82[30:0];
  assign GEN_9 = {{1'd0}, T_88};
  assign T_89 = GEN_9 << 1;
  assign T_91 = T_89 & 32'haaaaaaaa;
  assign T_92 = T_87 | T_91;
  assign shin = T_41 ? io_in1 : T_92;
  assign T_94 = shin[31];
  assign T_95 = T_15 & T_94;
  assign T_96 = {T_95,shin};
  assign T_97 = $signed(T_96);
  assign T_98 = ($signed(T_97) >>> shamt) ;//($signed(T_97) >> shamt) | ; //$signed(T_97) >>> shamt;//$signed(T_97) >>> shamt;
  assign shout_r = T_98[31:0];
  assign T_103 = shout_r[31:16];
  assign T_104 = {{16'd0}, T_103};
  assign T_105 = shout_r[15:0];
  assign GEN_10 = {{16'd0}, T_105};
  assign T_106 = GEN_10 << 16;
  assign T_108 = T_106 & 32'hffff0000;
  assign T_109 = T_104 | T_108;
  assign T_113 = T_109[31:8];
  assign GEN_11 = {{8'd0}, T_113};
  assign T_114 = GEN_11 & 32'hff00ff;
  assign T_115 = T_109[23:0];
  assign GEN_12 = {{8'd0}, T_115};
  assign T_116 = GEN_12 << 8;
  assign T_118 = T_116 & 32'hff00ff00;
  assign T_119 = T_114 | T_118;
  assign T_123 = T_119[31:4];
  assign GEN_13 = {{4'd0}, T_123};
  assign T_124 = GEN_13 & 32'hf0f0f0f;
  assign T_125 = T_119[27:0];
  assign GEN_14 = {{4'd0}, T_125};
  assign T_126 = GEN_14 << 4;
  assign T_128 = T_126 & 32'hf0f0f0f0;
  assign T_129 = T_124 | T_128;
  assign T_133 = T_129[31:2];
  assign GEN_15 = {{2'd0}, T_133};
  assign T_134 = GEN_15 & 32'h33333333;
  assign T_135 = T_129[29:0];
  assign GEN_16 = {{2'd0}, T_135};
  assign T_136 = GEN_16 << 2;
  assign T_138 = T_136 & 32'hcccccccc;
  assign T_139 = T_134 | T_138;
  assign T_143 = T_139[31:1];
  assign GEN_17 = {{1'd0}, T_143};
  assign T_144 = GEN_17 & 32'h55555555;
  assign T_145 = T_139[30:0];
  assign GEN_18 = {{1'd0}, T_145};
  assign T_146 = GEN_18 << 1;
  assign T_148 = T_146 & 32'haaaaaaaa;
  assign shout_l = T_144 | T_148;
  assign T_153 = T_41 ? shout_r : 32'h0;
  assign T_154 = io_fn == 4'h1;
  assign T_156 = T_154 ? shout_l : 32'h0;
  assign shout = T_153 | T_156;
  assign T_157 = io_fn == 4'h4;
  assign T_158 = io_fn == 4'h6;
  assign T_159 = T_157 | T_158;
  assign T_161 = T_159 ? in1_xor_in2 : 32'h0;
  assign T_163 = io_fn == 4'h7;
  assign T_164 = T_158 | T_163;
  assign T_165 = io_in1 & io_in2;
  assign T_167 = T_164 ? T_165 : 32'h0;
  assign logic$ = T_161 | T_167;
  assign T_168 = io_fn == 4'h2;
  assign T_169 = io_fn == 4'h3;
  assign T_170 = T_168 | T_169;
  assign T_171 = io_fn >= 4'hc;
  assign T_172 = T_170 | T_171;
  assign T_173 = T_172 & io_cmp_out;
  assign GEN_19 = {{31'd0}, T_173};
  assign T_174 = GEN_19 | logic$;
  assign shift_logic = T_174 | shout;
  assign T_175 = io_fn == 4'h0;
  assign T_176 = io_fn == 4'ha;
  assign T_177 = T_175 | T_176;
  assign out = T_177 ? io_adder_out : shift_logic;
endmodule