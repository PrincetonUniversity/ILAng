module GB(
arg_0_TREADY,
arg_1_TDATA,
arg_1_TVALID,
LB1D_buff,
LB1D_p_cnt,
LB2D_proc_w,
LB2D_proc_x,
LB2D_proc_y,
LB2D_shift_0,
LB2D_shift_1,
LB2D_shift_2,
LB2D_shift_3,
LB2D_shift_4,
LB2D_shift_5,
LB2D_shift_6,
LB2D_shift_7,
LB2D_shift_x,
LB2D_shift_y,
arg_0_TDATA,
arg_0_TVALID,
arg_1_TREADY,
gb_exit_it_1,
gb_exit_it_2,
gb_exit_it_3,
gb_exit_it_4,
gb_exit_it_5,
gb_exit_it_6,
gb_exit_it_7,
gb_exit_it_8,
gb_p_cnt,
gb_pp_it_1,
gb_pp_it_2,
gb_pp_it_3,
gb_pp_it_4,
gb_pp_it_5,
gb_pp_it_6,
gb_pp_it_7,
gb_pp_it_8,
gb_pp_it_9,
in_stream_buff_0,
in_stream_buff_1,
in_stream_empty,
in_stream_full,
slice_stream_buff_0,
slice_stream_buff_1,
slice_stream_empty,
slice_stream_full,
stencil_stream_buff_0,
stencil_stream_buff_1,
stencil_stream_empty,
stencil_stream_full,
clk,rst,
step
);
input            arg_0_TREADY;
input      [7:0] arg_1_TDATA;
input            arg_1_TVALID;
input clk;
input rst;
input step;
output      [7:0] LB1D_buff;
output     [18:0] LB1D_p_cnt;
output     [63:0] LB2D_proc_w;
output      [8:0] LB2D_proc_x;
output      [9:0] LB2D_proc_y;
output     [71:0] LB2D_shift_0;
output     [71:0] LB2D_shift_1;
output     [71:0] LB2D_shift_2;
output     [71:0] LB2D_shift_3;
output     [71:0] LB2D_shift_4;
output     [71:0] LB2D_shift_5;
output     [71:0] LB2D_shift_6;
output     [71:0] LB2D_shift_7;
output      [8:0] LB2D_shift_x;
output      [9:0] LB2D_shift_y;
output      [7:0] arg_0_TDATA;
output            arg_0_TVALID;
output            arg_1_TREADY;
output            gb_exit_it_1;
output            gb_exit_it_2;
output            gb_exit_it_3;
output            gb_exit_it_4;
output            gb_exit_it_5;
output            gb_exit_it_6;
output            gb_exit_it_7;
output            gb_exit_it_8;
output     [18:0] gb_p_cnt;
output            gb_pp_it_1;
output            gb_pp_it_2;
output            gb_pp_it_3;
output            gb_pp_it_4;
output            gb_pp_it_5;
output            gb_pp_it_6;
output            gb_pp_it_7;
output            gb_pp_it_8;
output            gb_pp_it_9;
output      [7:0] in_stream_buff_0;
output      [7:0] in_stream_buff_1;
output            in_stream_empty;
output            in_stream_full;
output     [71:0] slice_stream_buff_0;
output     [71:0] slice_stream_buff_1;
output            slice_stream_empty;
output            slice_stream_full;
output    [647:0] stencil_stream_buff_0;
output    [647:0] stencil_stream_buff_1;
output            stencil_stream_empty;
output            stencil_stream_full;
reg      [7:0] LB1D_buff;
reg     [18:0] LB1D_p_cnt;
reg     [63:0] LB2D_proc_w;
reg      [8:0] LB2D_proc_x;
reg      [9:0] LB2D_proc_y;
reg     [71:0] LB2D_shift_0;
reg     [71:0] LB2D_shift_1;
reg     [71:0] LB2D_shift_2;
reg     [71:0] LB2D_shift_3;
reg     [71:0] LB2D_shift_4;
reg     [71:0] LB2D_shift_5;
reg     [71:0] LB2D_shift_6;
reg     [71:0] LB2D_shift_7;
reg      [8:0] LB2D_shift_x;
reg      [9:0] LB2D_shift_y;
reg      [7:0] arg_0_TDATA;
reg            arg_0_TVALID;
reg            arg_1_TREADY;
reg            gb_exit_it_1;
reg            gb_exit_it_2;
reg            gb_exit_it_3;
reg            gb_exit_it_4;
reg            gb_exit_it_5;
reg            gb_exit_it_6;
reg            gb_exit_it_7;
reg            gb_exit_it_8;
reg     [18:0] gb_p_cnt;
reg            gb_pp_it_1;
reg            gb_pp_it_2;
reg            gb_pp_it_3;
reg            gb_pp_it_4;
reg            gb_pp_it_5;
reg            gb_pp_it_6;
reg            gb_pp_it_7;
reg            gb_pp_it_8;
reg            gb_pp_it_9;
reg      [7:0] in_stream_buff_0;
reg      [7:0] in_stream_buff_1;
reg            in_stream_empty;
reg            in_stream_full;
reg     [71:0] slice_stream_buff_0;
reg     [71:0] slice_stream_buff_1;
reg            slice_stream_empty;
reg            slice_stream_full;
reg    [647:0] stencil_stream_buff_0;
reg    [647:0] stencil_stream_buff_1;
reg            stencil_stream_empty;
reg            stencil_stream_full;
wire            arg_0_TREADY;
wire      [7:0] arg_1_TDATA;
wire            arg_1_TVALID;
wire            n0;
wire            n1;
wire            n2;
wire            n3;
wire            n4;
wire            n5;
wire            n6;
wire            n7;
wire            n8;
wire            n9;
wire            n10;
wire            n11;
wire            n12;
wire            n13;
wire            n14;
wire            n15;
wire            n16;
wire            n17;
wire            n18;
wire            n19;
wire            n20;
wire            n21;
wire            n22;
wire            n23;
wire            n24;
wire            n25;
wire            n26;
wire            n27;
wire            n28;
wire            n29;
wire            n30;
wire            n31;
wire            n32;
wire            n33;
wire      [7:0] n34;
wire      [7:0] n35;
wire      [7:0] n36;
wire      [7:0] n37;
wire      [7:0] n38;
wire      [7:0] n39;
wire     [18:0] n40;
wire     [18:0] n41;
wire     [18:0] n42;
wire     [18:0] n43;
wire     [18:0] n44;
wire     [18:0] n45;
wire     [18:0] n46;
wire            n47;
wire            n48;
wire     [63:0] n49;
wire     [63:0] n50;
wire     [63:0] n51;
wire     [63:0] n52;
wire     [63:0] n53;
wire     [63:0] n54;
wire     [63:0] n55;
wire     [63:0] n56;
wire     [63:0] n57;
wire      [8:0] n58;
wire      [8:0] n59;
wire      [8:0] n60;
wire      [8:0] n61;
wire      [8:0] n62;
wire      [8:0] n63;
wire      [8:0] n64;
wire      [8:0] n65;
wire            n66;
wire      [9:0] n67;
wire      [9:0] n68;
wire      [9:0] n69;
wire      [9:0] n70;
wire      [9:0] n71;
wire      [9:0] n72;
wire      [9:0] n73;
wire      [9:0] n74;
wire      [9:0] n75;
wire            n76;
wire     [71:0] n77;
wire     [71:0] n78;
wire     [71:0] n79;
wire     [71:0] n80;
wire     [71:0] n81;
wire     [71:0] n82;
wire     [71:0] n83;
wire     [71:0] n84;
wire     [71:0] n85;
wire     [71:0] n86;
wire     [71:0] n87;
wire     [71:0] n88;
wire     [71:0] n89;
wire     [71:0] n90;
wire     [71:0] n91;
wire     [71:0] n92;
wire     [71:0] n93;
wire     [71:0] n94;
wire     [71:0] n95;
wire     [71:0] n96;
wire     [71:0] n97;
wire     [71:0] n98;
wire     [71:0] n99;
wire     [71:0] n100;
wire     [71:0] n101;
wire     [71:0] n102;
wire     [71:0] n103;
wire     [71:0] n104;
wire     [71:0] n105;
wire     [71:0] n106;
wire     [71:0] n107;
wire     [71:0] n108;
wire     [71:0] n109;
wire     [71:0] n110;
wire     [71:0] n111;
wire     [71:0] n112;
wire     [71:0] n113;
wire     [71:0] n114;
wire     [71:0] n115;
wire     [71:0] n116;
wire     [71:0] n117;
wire     [71:0] n118;
wire     [71:0] n119;
wire     [71:0] n120;
wire     [71:0] n121;
wire     [71:0] n122;
wire     [71:0] n123;
wire     [71:0] n124;
wire     [71:0] n125;
wire            n126;
wire      [8:0] n127;
wire      [8:0] n128;
wire      [8:0] n129;
wire      [8:0] n130;
wire      [8:0] n131;
wire      [8:0] n132;
wire      [8:0] n133;
wire      [8:0] n134;
wire            n135;
wire      [9:0] n136;
wire      [9:0] n137;
wire      [9:0] n138;
wire      [9:0] n139;
wire      [9:0] n140;
wire      [9:0] n141;
wire      [9:0] n142;
wire      [9:0] n143;
wire      [9:0] n144;
wire            n145;
wire    [647:0] n146;
wire      [7:0] n147;
wire      [7:0] n148;
wire      [7:0] n149;
wire      [7:0] n150;
wire      [7:0] n151;
wire      [7:0] n152;
wire      [7:0] n153;
wire            n154;
wire            n155;
wire            n156;
wire            n157;
wire            n158;
wire            n159;
wire            n160;
wire            n161;
wire            n162;
wire            n163;
wire            n164;
wire            n165;
wire            n166;
wire            n167;
wire     [18:0] n168;
wire            n169;
wire            n170;
wire            n171;
wire            n172;
wire            n173;
wire            n174;
wire            n175;
wire            n176;
wire            n177;
wire            n178;
wire            n179;
wire            n180;
wire            n181;
wire            n182;
wire            n183;
wire            n184;
wire            n185;
wire            n186;
wire            n187;
wire            n188;
wire            n189;
wire            n190;
wire            n191;
wire            n192;
wire            n193;
wire            n194;
wire            n195;
wire            n196;
wire            n197;
wire            n198;
wire            n199;
wire            n200;
wire            n201;
wire            n202;
wire            n203;
wire            n204;
wire            n205;
wire            n206;
wire            n207;
wire            n208;
wire            n209;
wire            n210;
wire            n211;
wire            n212;
wire            n213;
wire            n214;
wire            n215;
wire            n216;
wire            n217;
wire            n218;
wire            n219;
wire     [18:0] n220;
wire     [18:0] n221;
wire     [18:0] n222;
wire     [18:0] n223;
wire     [18:0] n224;
wire     [18:0] n225;
wire     [18:0] n226;
wire            n227;
wire            n228;
wire            n229;
wire            n230;
wire            n231;
wire            n232;
wire            n233;
wire            n234;
wire            n235;
wire            n236;
wire            n237;
wire            n238;
wire            n239;
wire            n240;
wire            n241;
wire            n242;
wire            n243;
wire            n244;
wire            n245;
wire            n246;
wire            n247;
wire            n248;
wire            n249;
wire            n250;
wire            n251;
wire            n252;
wire            n253;
wire            n254;
wire            n255;
wire            n256;
wire            n257;
wire            n258;
wire            n259;
wire            n260;
wire            n261;
wire            n262;
wire            n263;
wire            n264;
wire            n265;
wire            n266;
wire            n267;
wire            n268;
wire            n269;
wire            n270;
wire            n271;
wire            n272;
wire            n273;
wire            n274;
wire            n275;
wire            n276;
wire            n277;
wire            n278;
wire            n279;
wire            n280;
wire      [7:0] n281;
wire      [7:0] n282;
wire      [7:0] n283;
wire      [7:0] n284;
wire      [7:0] n285;
wire      [7:0] n286;
wire      [7:0] n287;
wire      [7:0] n288;
wire      [7:0] n289;
wire      [7:0] n290;
wire      [7:0] n291;
wire      [7:0] n292;
wire            n293;
wire            n294;
wire            n295;
wire            n296;
wire            n297;
wire            n298;
wire            n299;
wire            n300;
wire            n301;
wire            n302;
wire            n303;
wire            n304;
wire            n305;
wire            n306;
wire            n307;
wire            n308;
wire      [7:0] n309;
wire            n310;
wire      [7:0] n311;
wire            n312;
wire      [7:0] n313;
wire            n314;
wire      [7:0] n315;
wire            n316;
wire      [7:0] n317;
wire            n318;
wire      [7:0] n319;
wire            n320;
wire      [7:0] n321;
wire            n322;
wire      [7:0] n323;
wire      [7:0] n324;
wire      [7:0] n325;
wire      [7:0] n326;
wire      [7:0] n327;
wire      [7:0] n328;
wire      [7:0] n329;
wire      [7:0] n330;
wire      [7:0] n331;
wire      [7:0] n332;
wire      [7:0] n333;
wire      [7:0] n334;
wire      [7:0] n335;
wire      [7:0] n336;
wire      [7:0] n337;
wire      [7:0] n338;
wire      [7:0] n339;
wire      [7:0] n340;
wire      [7:0] n341;
wire      [7:0] n342;
wire      [7:0] n343;
wire      [7:0] n344;
wire      [7:0] n345;
wire      [7:0] n346;
wire      [7:0] n347;
wire      [7:0] n348;
wire      [7:0] n349;
wire      [7:0] n350;
wire      [7:0] n351;
wire      [7:0] n352;
wire      [7:0] n353;
wire      [7:0] n354;
wire      [7:0] n355;
wire      [7:0] n356;
wire      [7:0] n357;
wire      [7:0] n358;
wire      [7:0] n359;
wire      [7:0] n360;
wire      [7:0] n361;
wire      [7:0] n362;
wire      [7:0] n363;
wire      [7:0] n364;
wire      [7:0] n365;
wire      [7:0] n366;
wire      [7:0] n367;
wire      [7:0] n368;
wire      [7:0] n369;
wire      [7:0] n370;
wire      [7:0] n371;
wire      [7:0] n372;
wire      [7:0] n373;
wire      [7:0] n374;
wire      [7:0] n375;
wire      [7:0] n376;
wire      [7:0] n377;
wire      [7:0] n378;
wire      [7:0] n379;
wire      [7:0] n380;
wire     [15:0] n381;
wire     [23:0] n382;
wire     [31:0] n383;
wire     [39:0] n384;
wire     [47:0] n385;
wire     [55:0] n386;
wire     [63:0] n387;
wire     [71:0] n388;
wire     [71:0] n389;
wire     [71:0] n390;
wire     [71:0] n391;
wire     [71:0] n392;
wire     [71:0] n393;
wire     [71:0] n394;
wire     [71:0] n395;
wire     [71:0] n396;
wire     [71:0] n397;
wire     [71:0] n398;
wire     [71:0] n399;
wire     [71:0] n400;
wire     [71:0] n401;
wire     [71:0] n402;
wire            n403;
wire            n404;
wire            n405;
wire            n406;
wire            n407;
wire            n408;
wire            n409;
wire            n410;
wire            n411;
wire            n412;
wire            n413;
wire            n414;
wire            n415;
wire            n416;
wire            n417;
wire            n418;
wire            n419;
wire            n420;
wire      [7:0] n421;
wire      [7:0] n422;
wire      [7:0] n423;
wire      [7:0] n424;
wire      [7:0] n425;
wire      [7:0] n426;
wire      [7:0] n427;
wire      [7:0] n428;
wire      [7:0] n429;
wire     [15:0] n430;
wire     [23:0] n431;
wire     [31:0] n432;
wire     [39:0] n433;
wire     [47:0] n434;
wire     [55:0] n435;
wire     [63:0] n436;
wire     [71:0] n437;
wire      [7:0] n438;
wire      [7:0] n439;
wire      [7:0] n440;
wire      [7:0] n441;
wire      [7:0] n442;
wire      [7:0] n443;
wire      [7:0] n444;
wire      [7:0] n445;
wire      [7:0] n446;
wire     [15:0] n447;
wire     [23:0] n448;
wire     [31:0] n449;
wire     [39:0] n450;
wire     [47:0] n451;
wire     [55:0] n452;
wire     [63:0] n453;
wire     [71:0] n454;
wire      [7:0] n455;
wire      [7:0] n456;
wire      [7:0] n457;
wire      [7:0] n458;
wire      [7:0] n459;
wire      [7:0] n460;
wire      [7:0] n461;
wire      [7:0] n462;
wire      [7:0] n463;
wire     [15:0] n464;
wire     [23:0] n465;
wire     [31:0] n466;
wire     [39:0] n467;
wire     [47:0] n468;
wire     [55:0] n469;
wire     [63:0] n470;
wire     [71:0] n471;
wire      [7:0] n472;
wire      [7:0] n473;
wire      [7:0] n474;
wire      [7:0] n475;
wire      [7:0] n476;
wire      [7:0] n477;
wire      [7:0] n478;
wire      [7:0] n479;
wire      [7:0] n480;
wire     [15:0] n481;
wire     [23:0] n482;
wire     [31:0] n483;
wire     [39:0] n484;
wire     [47:0] n485;
wire     [55:0] n486;
wire     [63:0] n487;
wire     [71:0] n488;
wire      [7:0] n489;
wire      [7:0] n490;
wire      [7:0] n491;
wire      [7:0] n492;
wire      [7:0] n493;
wire      [7:0] n494;
wire      [7:0] n495;
wire      [7:0] n496;
wire      [7:0] n497;
wire     [15:0] n498;
wire     [23:0] n499;
wire     [31:0] n500;
wire     [39:0] n501;
wire     [47:0] n502;
wire     [55:0] n503;
wire     [63:0] n504;
wire     [71:0] n505;
wire      [7:0] n506;
wire      [7:0] n507;
wire      [7:0] n508;
wire      [7:0] n509;
wire      [7:0] n510;
wire      [7:0] n511;
wire      [7:0] n512;
wire      [7:0] n513;
wire      [7:0] n514;
wire     [15:0] n515;
wire     [23:0] n516;
wire     [31:0] n517;
wire     [39:0] n518;
wire     [47:0] n519;
wire     [55:0] n520;
wire     [63:0] n521;
wire     [71:0] n522;
wire      [7:0] n523;
wire      [7:0] n524;
wire      [7:0] n525;
wire      [7:0] n526;
wire      [7:0] n527;
wire      [7:0] n528;
wire      [7:0] n529;
wire      [7:0] n530;
wire      [7:0] n531;
wire     [15:0] n532;
wire     [23:0] n533;
wire     [31:0] n534;
wire     [39:0] n535;
wire     [47:0] n536;
wire     [55:0] n537;
wire     [63:0] n538;
wire     [71:0] n539;
wire      [7:0] n540;
wire      [7:0] n541;
wire      [7:0] n542;
wire      [7:0] n543;
wire      [7:0] n544;
wire      [7:0] n545;
wire      [7:0] n546;
wire      [7:0] n547;
wire      [7:0] n548;
wire     [15:0] n549;
wire     [23:0] n550;
wire     [31:0] n551;
wire     [39:0] n552;
wire     [47:0] n553;
wire     [55:0] n554;
wire     [63:0] n555;
wire     [71:0] n556;
wire      [7:0] n557;
wire      [7:0] n558;
wire      [7:0] n559;
wire      [7:0] n560;
wire      [7:0] n561;
wire      [7:0] n562;
wire      [7:0] n563;
wire      [7:0] n564;
wire      [7:0] n565;
wire     [15:0] n566;
wire     [23:0] n567;
wire     [31:0] n568;
wire     [39:0] n569;
wire     [47:0] n570;
wire     [55:0] n571;
wire     [63:0] n572;
wire     [71:0] n573;
wire    [143:0] n574;
wire    [215:0] n575;
wire    [287:0] n576;
wire    [359:0] n577;
wire    [431:0] n578;
wire    [503:0] n579;
wire    [575:0] n580;
wire    [647:0] n581;
wire    [647:0] n582;
wire    [647:0] n583;
wire    [647:0] n584;
wire    [647:0] n585;
wire    [647:0] n586;
wire    [647:0] n587;
wire    [647:0] n588;
wire    [647:0] n589;
wire    [647:0] n590;
wire    [647:0] n591;
wire    [647:0] n592;
wire    [647:0] n593;
wire    [647:0] n594;
wire            n595;
wire            n596;
wire            n597;
wire            n598;
wire            n599;
wire            n600;
wire            n601;
wire            n602;
wire            n603;
wire            n604;
wire            n605;
wire            n606;
wire            n607;
wire            n608;
wire            n609;
wire            n610;
wire            n611;
wire            n612;
wire      [8:0] LB2D_proc_0_addr0;
wire      [7:0] LB2D_proc_0_data0;
wire            n613;
wire            n614;
wire            n615;
wire            n616;
wire            n617;
wire            n618;
wire            n619;
wire            n620;
wire            n621;
wire            n622;
wire            n623;
wire            n624;
wire            n625;
wire            n626;
wire            n627;
wire            n628;
wire            n629;
wire            n630;
wire            n631;
wire      [8:0] LB2D_proc_1_addr0;
wire      [7:0] LB2D_proc_1_data0;
wire            n632;
wire            n633;
wire            n634;
wire      [8:0] LB2D_proc_2_addr0;
wire      [7:0] LB2D_proc_2_data0;
wire            n635;
wire            n636;
wire            n637;
wire      [8:0] LB2D_proc_3_addr0;
wire      [7:0] LB2D_proc_3_data0;
wire            n638;
wire            n639;
wire            n640;
wire      [8:0] LB2D_proc_4_addr0;
wire      [7:0] LB2D_proc_4_data0;
wire            n641;
wire            n642;
wire            n643;
wire      [8:0] LB2D_proc_5_addr0;
wire      [7:0] LB2D_proc_5_data0;
wire            n644;
wire            n645;
wire            n646;
wire      [8:0] LB2D_proc_6_addr0;
wire      [7:0] LB2D_proc_6_data0;
wire            n647;
wire            n648;
wire            n649;
wire      [8:0] LB2D_proc_7_addr0;
wire      [7:0] LB2D_proc_7_data0;
wire            n650;
wire            n651;
wire            n652;
wire            n653;
reg      [7:0] LB2D_proc_0[511:0];
reg      [7:0] LB2D_proc_1[511:0];
reg      [7:0] LB2D_proc_2[511:0];
reg      [7:0] LB2D_proc_3[511:0];
reg      [7:0] LB2D_proc_4[511:0];
reg      [7:0] LB2D_proc_5[511:0];
reg      [7:0] LB2D_proc_6[511:0];
reg      [7:0] LB2D_proc_7[511:0];
wire clk;
wire rst;
wire step;
assign n0 =  ( arg_0_TREADY ) == ( 1'd1 )  ;
assign n1 =  ( arg_0_TVALID ) == ( 1'd1 )  ;
assign n2 =  ( n0 ) & ( n1 )  ;
assign n3 =  ( arg_1_TVALID ) == ( 1'd0 )  ;
assign n4 =  ( n2 ) & ( n3 )  ;
assign n5 =  ( arg_1_TREADY ) == ( 1'd1 )  ;
assign n6 =  ( arg_1_TVALID ) == ( 1'd1 )  ;
assign n7 =  ( n5 ) & ( n6 )  ;
assign n8 =  ( arg_0_TREADY ) == ( 1'd0 )  ;
assign n9 =  ( n7 ) & ( n8 )  ;
assign n10 =  ( arg_0_TVALID ) == ( 1'd0 )  ;
assign n11 =  ( gb_exit_it_1 ) == ( 1'd0 )  ;
assign n12 =  ( stencil_stream_empty ) == ( 1'd0 )  ;
assign n13 =  ( n11 ) & ( n12 )  ;
assign n14 =  ( gb_exit_it_1 ) == ( 1'd1 )  ;
assign n15 =  ( gb_exit_it_8 ) == ( 1'd0 )  ;
assign n16 =  ( n14 ) & ( n15 )  ;
assign n17 =  ( n13 ) | ( n16 )  ;
assign n18 =  ( n10 ) & ( n17 )  ;
assign n19 =  ( slice_stream_empty ) == ( 1'd0 )  ;
assign n20 =  ( stencil_stream_full ) == ( 1'd0 )  ;
assign n21 =  ( LB2D_shift_x ) < ( 9'd8 )  ;
assign n22 =  ( n20 ) | ( n21 )  ;
assign n23 =  ( n19 ) & ( n22 )  ;
assign n24 =  ( in_stream_empty ) == ( 1'd0 )  ;
assign n25 =  ( slice_stream_full ) == ( 1'd0 )  ;
assign n26 =  ( LB2D_proc_y ) < ( 10'd8 )  ;
assign n27 =  ( n25 ) | ( n26 )  ;
assign n28 =  ( n24 ) & ( n27 )  ;
assign n29 =  ( arg_1_TREADY ) == ( 1'd0 )  ;
assign n30 =  ( in_stream_full ) == ( 1'd0 )  ;
assign n31 =  ( n29 ) & ( n30 )  ;
assign n32 =  ( LB1D_p_cnt ) != ( 19'd316224 )  ;
assign n33 =  ( n31 ) & ( n32 )  ;
assign n34 =  ( n33 ) ? ( LB1D_buff ) : ( LB1D_buff ) ;
assign n35 =  ( n28 ) ? ( LB1D_buff ) : ( n34 ) ;
assign n36 =  ( n23 ) ? ( LB1D_buff ) : ( n35 ) ;
assign n37 =  ( n18 ) ? ( LB1D_buff ) : ( n36 ) ;
assign n38 =  ( n9 ) ? ( arg_1_TDATA ) : ( n37 ) ;
assign n39 =  ( n4 ) ? ( arg_1_TDATA ) : ( n38 ) ;
assign n40 =  ( LB1D_p_cnt ) + ( 19'd1 )  ;
assign n41 =  ( n33 ) ? ( n40 ) : ( LB1D_p_cnt ) ;
assign n42 =  ( n28 ) ? ( LB1D_p_cnt ) : ( n41 ) ;
assign n43 =  ( n23 ) ? ( LB1D_p_cnt ) : ( n42 ) ;
assign n44 =  ( n18 ) ? ( LB1D_p_cnt ) : ( n43 ) ;
assign n45 =  ( n9 ) ? ( LB1D_p_cnt ) : ( n44 ) ;
assign n46 =  ( n4 ) ? ( LB1D_p_cnt ) : ( n45 ) ;
assign n47 =  ( LB2D_proc_w ) < ( 64'd7 )  ;
assign n48 =  ( LB2D_proc_x ) < ( 9'd487 )  ;
assign n49 =  ( LB2D_proc_w ) + ( 64'd1 )  ;
assign n50 =  ( n48 ) ? ( LB2D_proc_w ) : ( n49 ) ;
assign n51 =  ( n47 ) ? ( n50 ) : ( 64'd0 ) ;
assign n52 =  ( n33 ) ? ( LB2D_proc_w ) : ( LB2D_proc_w ) ;
assign n53 =  ( n28 ) ? ( n51 ) : ( n52 ) ;
assign n54 =  ( n23 ) ? ( LB2D_proc_w ) : ( n53 ) ;
assign n55 =  ( n18 ) ? ( LB2D_proc_w ) : ( n54 ) ;
assign n56 =  ( n9 ) ? ( LB2D_proc_w ) : ( n55 ) ;
assign n57 =  ( n4 ) ? ( LB2D_proc_w ) : ( n56 ) ;
assign n58 =  ( LB2D_proc_x ) + ( 9'd1 )  ;
assign n59 =  ( n48 ) ? ( n58 ) : ( 9'd0 ) ;
assign n60 =  ( n33 ) ? ( LB2D_proc_x ) : ( LB2D_proc_x ) ;
assign n61 =  ( n28 ) ? ( n59 ) : ( n60 ) ;
assign n62 =  ( n23 ) ? ( LB2D_proc_x ) : ( n61 ) ;
assign n63 =  ( n18 ) ? ( LB2D_proc_x ) : ( n62 ) ;
assign n64 =  ( n9 ) ? ( LB2D_proc_x ) : ( n63 ) ;
assign n65 =  ( n4 ) ? ( LB2D_proc_x ) : ( n64 ) ;
assign n66 =  ( LB2D_proc_y ) < ( 10'd487 )  ;
assign n67 =  ( LB2D_proc_y ) + ( 10'd1 )  ;
assign n68 =  ( n48 ) ? ( LB2D_proc_y ) : ( n67 ) ;
assign n69 =  ( n66 ) ? ( n68 ) : ( 10'd487 ) ;
assign n70 =  ( n33 ) ? ( LB2D_proc_y ) : ( LB2D_proc_y ) ;
assign n71 =  ( n28 ) ? ( n69 ) : ( n70 ) ;
assign n72 =  ( n23 ) ? ( LB2D_proc_y ) : ( n71 ) ;
assign n73 =  ( n18 ) ? ( LB2D_proc_y ) : ( n72 ) ;
assign n74 =  ( n9 ) ? ( LB2D_proc_y ) : ( n73 ) ;
assign n75 =  ( n4 ) ? ( LB2D_proc_y ) : ( n74 ) ;
assign n76 =  ( slice_stream_full ) == ( 1'd1 )  ;
assign n77 =  ( n76 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n78 =  ( n33 ) ? ( LB2D_shift_0 ) : ( LB2D_shift_0 ) ;
assign n79 =  ( n28 ) ? ( LB2D_shift_0 ) : ( n78 ) ;
assign n80 =  ( n23 ) ? ( n77 ) : ( n79 ) ;
assign n81 =  ( n18 ) ? ( LB2D_shift_0 ) : ( n80 ) ;
assign n82 =  ( n9 ) ? ( LB2D_shift_0 ) : ( n81 ) ;
assign n83 =  ( n4 ) ? ( LB2D_shift_0 ) : ( n82 ) ;
assign n84 =  ( n33 ) ? ( LB2D_shift_1 ) : ( LB2D_shift_1 ) ;
assign n85 =  ( n28 ) ? ( LB2D_shift_1 ) : ( n84 ) ;
assign n86 =  ( n23 ) ? ( LB2D_shift_0 ) : ( n85 ) ;
assign n87 =  ( n18 ) ? ( LB2D_shift_1 ) : ( n86 ) ;
assign n88 =  ( n9 ) ? ( LB2D_shift_1 ) : ( n87 ) ;
assign n89 =  ( n4 ) ? ( LB2D_shift_1 ) : ( n88 ) ;
assign n90 =  ( n33 ) ? ( LB2D_shift_2 ) : ( LB2D_shift_2 ) ;
assign n91 =  ( n28 ) ? ( LB2D_shift_2 ) : ( n90 ) ;
assign n92 =  ( n23 ) ? ( LB2D_shift_1 ) : ( n91 ) ;
assign n93 =  ( n18 ) ? ( LB2D_shift_2 ) : ( n92 ) ;
assign n94 =  ( n9 ) ? ( LB2D_shift_2 ) : ( n93 ) ;
assign n95 =  ( n4 ) ? ( LB2D_shift_2 ) : ( n94 ) ;
assign n96 =  ( n33 ) ? ( LB2D_shift_3 ) : ( LB2D_shift_3 ) ;
assign n97 =  ( n28 ) ? ( LB2D_shift_3 ) : ( n96 ) ;
assign n98 =  ( n23 ) ? ( LB2D_shift_2 ) : ( n97 ) ;
assign n99 =  ( n18 ) ? ( LB2D_shift_3 ) : ( n98 ) ;
assign n100 =  ( n9 ) ? ( LB2D_shift_3 ) : ( n99 ) ;
assign n101 =  ( n4 ) ? ( LB2D_shift_3 ) : ( n100 ) ;
assign n102 =  ( n33 ) ? ( LB2D_shift_4 ) : ( LB2D_shift_4 ) ;
assign n103 =  ( n28 ) ? ( LB2D_shift_4 ) : ( n102 ) ;
assign n104 =  ( n23 ) ? ( LB2D_shift_3 ) : ( n103 ) ;
assign n105 =  ( n18 ) ? ( LB2D_shift_4 ) : ( n104 ) ;
assign n106 =  ( n9 ) ? ( LB2D_shift_4 ) : ( n105 ) ;
assign n107 =  ( n4 ) ? ( LB2D_shift_4 ) : ( n106 ) ;
assign n108 =  ( n33 ) ? ( LB2D_shift_5 ) : ( LB2D_shift_5 ) ;
assign n109 =  ( n28 ) ? ( LB2D_shift_5 ) : ( n108 ) ;
assign n110 =  ( n23 ) ? ( LB2D_shift_4 ) : ( n109 ) ;
assign n111 =  ( n18 ) ? ( LB2D_shift_5 ) : ( n110 ) ;
assign n112 =  ( n9 ) ? ( LB2D_shift_5 ) : ( n111 ) ;
assign n113 =  ( n4 ) ? ( LB2D_shift_5 ) : ( n112 ) ;
assign n114 =  ( n33 ) ? ( LB2D_shift_6 ) : ( LB2D_shift_6 ) ;
assign n115 =  ( n28 ) ? ( LB2D_shift_6 ) : ( n114 ) ;
assign n116 =  ( n23 ) ? ( LB2D_shift_5 ) : ( n115 ) ;
assign n117 =  ( n18 ) ? ( LB2D_shift_6 ) : ( n116 ) ;
assign n118 =  ( n9 ) ? ( LB2D_shift_6 ) : ( n117 ) ;
assign n119 =  ( n4 ) ? ( LB2D_shift_6 ) : ( n118 ) ;
assign n120 =  ( n33 ) ? ( LB2D_shift_7 ) : ( LB2D_shift_7 ) ;
assign n121 =  ( n28 ) ? ( LB2D_shift_7 ) : ( n120 ) ;
assign n122 =  ( n23 ) ? ( LB2D_shift_6 ) : ( n121 ) ;
assign n123 =  ( n18 ) ? ( LB2D_shift_7 ) : ( n122 ) ;
assign n124 =  ( n9 ) ? ( LB2D_shift_7 ) : ( n123 ) ;
assign n125 =  ( n4 ) ? ( LB2D_shift_7 ) : ( n124 ) ;
assign n126 =  ( LB2D_shift_x ) < ( 9'd487 )  ;
assign n127 =  ( LB2D_shift_x ) + ( 9'd1 )  ;
assign n128 =  ( n126 ) ? ( n127 ) : ( 9'd0 ) ;
assign n129 =  ( n33 ) ? ( LB2D_shift_x ) : ( LB2D_shift_x ) ;
assign n130 =  ( n28 ) ? ( LB2D_shift_x ) : ( n129 ) ;
assign n131 =  ( n23 ) ? ( n128 ) : ( n130 ) ;
assign n132 =  ( n18 ) ? ( LB2D_shift_x ) : ( n131 ) ;
assign n133 =  ( n9 ) ? ( LB2D_shift_x ) : ( n132 ) ;
assign n134 =  ( n4 ) ? ( LB2D_shift_x ) : ( n133 ) ;
assign n135 =  ( LB2D_shift_y ) < ( 10'd479 )  ;
assign n136 =  ( LB2D_shift_y ) + ( 10'd1 )  ;
assign n137 =  ( n126 ) ? ( LB2D_shift_y ) : ( n136 ) ;
assign n138 =  ( n135 ) ? ( n137 ) : ( 10'd479 ) ;
assign n139 =  ( n33 ) ? ( LB2D_shift_y ) : ( LB2D_shift_y ) ;
assign n140 =  ( n28 ) ? ( LB2D_shift_y ) : ( n139 ) ;
assign n141 =  ( n23 ) ? ( n138 ) : ( n140 ) ;
assign n142 =  ( n18 ) ? ( LB2D_shift_y ) : ( n141 ) ;
assign n143 =  ( n9 ) ? ( LB2D_shift_y ) : ( n142 ) ;
assign n144 =  ( n4 ) ? ( LB2D_shift_y ) : ( n143 ) ;
assign n145 =  ( stencil_stream_full ) == ( 1'd1 )  ;
assign n146 =  ( n145 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_0 ) ;
//assign n147 = gb_fun(n146) ;
gb_fun gb_fun_U (
    .stencil (n146),
    .result (n147)
);

assign n148 =  ( n33 ) ? ( arg_0_TDATA ) : ( arg_0_TDATA ) ;
assign n149 =  ( n28 ) ? ( arg_0_TDATA ) : ( n148 ) ;
assign n150 =  ( n23 ) ? ( arg_0_TDATA ) : ( n149 ) ;
assign n151 =  ( n18 ) ? ( n147 ) : ( n150 ) ;
assign n152 =  ( n9 ) ? ( arg_0_TDATA ) : ( n151 ) ;
assign n153 =  ( n4 ) ? ( arg_0_TDATA ) : ( n152 ) ;
assign n154 =  ( gb_pp_it_8 ) == ( 1'd1 )  ;
assign n155 =  ( n154 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n156 =  ( n33 ) ? ( arg_0_TVALID ) : ( arg_0_TVALID ) ;
assign n157 =  ( n28 ) ? ( arg_0_TVALID ) : ( n156 ) ;
assign n158 =  ( n23 ) ? ( arg_0_TVALID ) : ( n157 ) ;
assign n159 =  ( n18 ) ? ( n155 ) : ( n158 ) ;
assign n160 =  ( n9 ) ? ( arg_0_TVALID ) : ( n159 ) ;
assign n161 =  ( n4 ) ? ( 1'd0 ) : ( n160 ) ;
assign n162 =  ( n33 ) ? ( 1'd1 ) : ( arg_1_TREADY ) ;
assign n163 =  ( n28 ) ? ( arg_1_TREADY ) : ( n162 ) ;
assign n164 =  ( n23 ) ? ( arg_1_TREADY ) : ( n163 ) ;
assign n165 =  ( n18 ) ? ( arg_1_TREADY ) : ( n164 ) ;
assign n166 =  ( n9 ) ? ( 1'd0 ) : ( n165 ) ;
assign n167 =  ( n4 ) ? ( 1'd0 ) : ( n166 ) ;
assign n168 =  ( gb_p_cnt ) + ( 19'd1 )  ;
assign n169 =  ( n168 ) == ( 19'd307200 )  ;
assign n170 =  ( n169 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n171 =  ( n33 ) ? ( gb_exit_it_1 ) : ( gb_exit_it_1 ) ;
assign n172 =  ( n28 ) ? ( gb_exit_it_1 ) : ( n171 ) ;
assign n173 =  ( n23 ) ? ( gb_exit_it_1 ) : ( n172 ) ;
assign n174 =  ( n18 ) ? ( n170 ) : ( n173 ) ;
assign n175 =  ( n9 ) ? ( gb_exit_it_1 ) : ( n174 ) ;
assign n176 =  ( n4 ) ? ( gb_exit_it_1 ) : ( n175 ) ;
assign n177 =  ( n33 ) ? ( gb_exit_it_2 ) : ( gb_exit_it_2 ) ;
assign n178 =  ( n28 ) ? ( gb_exit_it_2 ) : ( n177 ) ;
assign n179 =  ( n23 ) ? ( gb_exit_it_2 ) : ( n178 ) ;
assign n180 =  ( n18 ) ? ( gb_exit_it_1 ) : ( n179 ) ;
assign n181 =  ( n9 ) ? ( gb_exit_it_2 ) : ( n180 ) ;
assign n182 =  ( n4 ) ? ( gb_exit_it_2 ) : ( n181 ) ;
assign n183 =  ( n33 ) ? ( gb_exit_it_3 ) : ( gb_exit_it_3 ) ;
assign n184 =  ( n28 ) ? ( gb_exit_it_3 ) : ( n183 ) ;
assign n185 =  ( n23 ) ? ( gb_exit_it_3 ) : ( n184 ) ;
assign n186 =  ( n18 ) ? ( gb_exit_it_2 ) : ( n185 ) ;
assign n187 =  ( n9 ) ? ( gb_exit_it_3 ) : ( n186 ) ;
assign n188 =  ( n4 ) ? ( gb_exit_it_3 ) : ( n187 ) ;
assign n189 =  ( n33 ) ? ( gb_exit_it_4 ) : ( gb_exit_it_4 ) ;
assign n190 =  ( n28 ) ? ( gb_exit_it_4 ) : ( n189 ) ;
assign n191 =  ( n23 ) ? ( gb_exit_it_4 ) : ( n190 ) ;
assign n192 =  ( n18 ) ? ( gb_exit_it_3 ) : ( n191 ) ;
assign n193 =  ( n9 ) ? ( gb_exit_it_4 ) : ( n192 ) ;
assign n194 =  ( n4 ) ? ( gb_exit_it_4 ) : ( n193 ) ;
assign n195 =  ( n33 ) ? ( gb_exit_it_5 ) : ( gb_exit_it_5 ) ;
assign n196 =  ( n28 ) ? ( gb_exit_it_5 ) : ( n195 ) ;
assign n197 =  ( n23 ) ? ( gb_exit_it_5 ) : ( n196 ) ;
assign n198 =  ( n18 ) ? ( gb_exit_it_4 ) : ( n197 ) ;
assign n199 =  ( n9 ) ? ( gb_exit_it_5 ) : ( n198 ) ;
assign n200 =  ( n4 ) ? ( gb_exit_it_5 ) : ( n199 ) ;
assign n201 =  ( n33 ) ? ( gb_exit_it_6 ) : ( gb_exit_it_6 ) ;
assign n202 =  ( n28 ) ? ( gb_exit_it_6 ) : ( n201 ) ;
assign n203 =  ( n23 ) ? ( gb_exit_it_6 ) : ( n202 ) ;
assign n204 =  ( n18 ) ? ( gb_exit_it_5 ) : ( n203 ) ;
assign n205 =  ( n9 ) ? ( gb_exit_it_6 ) : ( n204 ) ;
assign n206 =  ( n4 ) ? ( gb_exit_it_6 ) : ( n205 ) ;
assign n207 =  ( n33 ) ? ( gb_exit_it_7 ) : ( gb_exit_it_7 ) ;
assign n208 =  ( n28 ) ? ( gb_exit_it_7 ) : ( n207 ) ;
assign n209 =  ( n23 ) ? ( gb_exit_it_7 ) : ( n208 ) ;
assign n210 =  ( n18 ) ? ( gb_exit_it_6 ) : ( n209 ) ;
assign n211 =  ( n9 ) ? ( gb_exit_it_7 ) : ( n210 ) ;
assign n212 =  ( n4 ) ? ( gb_exit_it_7 ) : ( n211 ) ;
assign n213 =  ( n33 ) ? ( gb_exit_it_8 ) : ( gb_exit_it_8 ) ;
assign n214 =  ( n28 ) ? ( gb_exit_it_8 ) : ( n213 ) ;
assign n215 =  ( n23 ) ? ( gb_exit_it_8 ) : ( n214 ) ;
assign n216 =  ( n18 ) ? ( gb_exit_it_7 ) : ( n215 ) ;
assign n217 =  ( n9 ) ? ( gb_exit_it_8 ) : ( n216 ) ;
assign n218 =  ( n4 ) ? ( gb_exit_it_8 ) : ( n217 ) ;
assign n219 =  ( gb_p_cnt ) < ( 19'd307200 )  ;
assign n220 =  ( n219 ) ? ( n168 ) : ( 19'd307200 ) ;
assign n221 =  ( n33 ) ? ( gb_p_cnt ) : ( gb_p_cnt ) ;
assign n222 =  ( n28 ) ? ( gb_p_cnt ) : ( n221 ) ;
assign n223 =  ( n23 ) ? ( gb_p_cnt ) : ( n222 ) ;
assign n224 =  ( n18 ) ? ( n220 ) : ( n223 ) ;
assign n225 =  ( n9 ) ? ( gb_p_cnt ) : ( n224 ) ;
assign n226 =  ( n4 ) ? ( gb_p_cnt ) : ( n225 ) ;
assign n227 =  ( n33 ) ? ( gb_pp_it_1 ) : ( gb_pp_it_1 ) ;
assign n228 =  ( n28 ) ? ( gb_pp_it_1 ) : ( n227 ) ;
assign n229 =  ( n23 ) ? ( gb_pp_it_1 ) : ( n228 ) ;
assign n230 =  ( n18 ) ? ( 1'd1 ) : ( n229 ) ;
assign n231 =  ( n9 ) ? ( gb_pp_it_1 ) : ( n230 ) ;
assign n232 =  ( n4 ) ? ( gb_pp_it_1 ) : ( n231 ) ;
assign n233 =  ( n33 ) ? ( gb_pp_it_2 ) : ( gb_pp_it_2 ) ;
assign n234 =  ( n28 ) ? ( gb_pp_it_2 ) : ( n233 ) ;
assign n235 =  ( n23 ) ? ( gb_pp_it_2 ) : ( n234 ) ;
assign n236 =  ( n18 ) ? ( gb_pp_it_1 ) : ( n235 ) ;
assign n237 =  ( n9 ) ? ( gb_pp_it_2 ) : ( n236 ) ;
assign n238 =  ( n4 ) ? ( gb_pp_it_2 ) : ( n237 ) ;
assign n239 =  ( n33 ) ? ( gb_pp_it_3 ) : ( gb_pp_it_3 ) ;
assign n240 =  ( n28 ) ? ( gb_pp_it_3 ) : ( n239 ) ;
assign n241 =  ( n23 ) ? ( gb_pp_it_3 ) : ( n240 ) ;
assign n242 =  ( n18 ) ? ( gb_pp_it_2 ) : ( n241 ) ;
assign n243 =  ( n9 ) ? ( gb_pp_it_3 ) : ( n242 ) ;
assign n244 =  ( n4 ) ? ( gb_pp_it_3 ) : ( n243 ) ;
assign n245 =  ( n33 ) ? ( gb_pp_it_4 ) : ( gb_pp_it_4 ) ;
assign n246 =  ( n28 ) ? ( gb_pp_it_4 ) : ( n245 ) ;
assign n247 =  ( n23 ) ? ( gb_pp_it_4 ) : ( n246 ) ;
assign n248 =  ( n18 ) ? ( gb_pp_it_3 ) : ( n247 ) ;
assign n249 =  ( n9 ) ? ( gb_pp_it_4 ) : ( n248 ) ;
assign n250 =  ( n4 ) ? ( gb_pp_it_4 ) : ( n249 ) ;
assign n251 =  ( n33 ) ? ( gb_pp_it_5 ) : ( gb_pp_it_5 ) ;
assign n252 =  ( n28 ) ? ( gb_pp_it_5 ) : ( n251 ) ;
assign n253 =  ( n23 ) ? ( gb_pp_it_5 ) : ( n252 ) ;
assign n254 =  ( n18 ) ? ( gb_pp_it_4 ) : ( n253 ) ;
assign n255 =  ( n9 ) ? ( gb_pp_it_5 ) : ( n254 ) ;
assign n256 =  ( n4 ) ? ( gb_pp_it_5 ) : ( n255 ) ;
assign n257 =  ( n33 ) ? ( gb_pp_it_6 ) : ( gb_pp_it_6 ) ;
assign n258 =  ( n28 ) ? ( gb_pp_it_6 ) : ( n257 ) ;
assign n259 =  ( n23 ) ? ( gb_pp_it_6 ) : ( n258 ) ;
assign n260 =  ( n18 ) ? ( gb_pp_it_5 ) : ( n259 ) ;
assign n261 =  ( n9 ) ? ( gb_pp_it_6 ) : ( n260 ) ;
assign n262 =  ( n4 ) ? ( gb_pp_it_6 ) : ( n261 ) ;
assign n263 =  ( n33 ) ? ( gb_pp_it_7 ) : ( gb_pp_it_7 ) ;
assign n264 =  ( n28 ) ? ( gb_pp_it_7 ) : ( n263 ) ;
assign n265 =  ( n23 ) ? ( gb_pp_it_7 ) : ( n264 ) ;
assign n266 =  ( n18 ) ? ( gb_pp_it_6 ) : ( n265 ) ;
assign n267 =  ( n9 ) ? ( gb_pp_it_7 ) : ( n266 ) ;
assign n268 =  ( n4 ) ? ( gb_pp_it_7 ) : ( n267 ) ;
assign n269 =  ( n33 ) ? ( gb_pp_it_8 ) : ( gb_pp_it_8 ) ;
assign n270 =  ( n28 ) ? ( gb_pp_it_8 ) : ( n269 ) ;
assign n271 =  ( n23 ) ? ( gb_pp_it_8 ) : ( n270 ) ;
assign n272 =  ( n18 ) ? ( gb_pp_it_7 ) : ( n271 ) ;
assign n273 =  ( n9 ) ? ( gb_pp_it_8 ) : ( n272 ) ;
assign n274 =  ( n4 ) ? ( gb_pp_it_8 ) : ( n273 ) ;
assign n275 =  ( n33 ) ? ( gb_pp_it_9 ) : ( gb_pp_it_9 ) ;
assign n276 =  ( n28 ) ? ( gb_pp_it_9 ) : ( n275 ) ;
assign n277 =  ( n23 ) ? ( gb_pp_it_9 ) : ( n276 ) ;
assign n278 =  ( n18 ) ? ( gb_pp_it_8 ) : ( n277 ) ;
assign n279 =  ( n9 ) ? ( gb_pp_it_9 ) : ( n278 ) ;
assign n280 =  ( n4 ) ? ( gb_pp_it_9 ) : ( n279 ) ;
assign n281 =  ( n33 ) ? ( LB1D_buff ) : ( in_stream_buff_0 ) ;
assign n282 =  ( n28 ) ? ( in_stream_buff_0 ) : ( n281 ) ;
assign n283 =  ( n23 ) ? ( in_stream_buff_0 ) : ( n282 ) ;
assign n284 =  ( n18 ) ? ( in_stream_buff_0 ) : ( n283 ) ;
assign n285 =  ( n9 ) ? ( in_stream_buff_0 ) : ( n284 ) ;
assign n286 =  ( n4 ) ? ( in_stream_buff_0 ) : ( n285 ) ;
assign n287 =  ( n33 ) ? ( in_stream_buff_0 ) : ( in_stream_buff_1 ) ;
assign n288 =  ( n28 ) ? ( in_stream_buff_1 ) : ( n287 ) ;
assign n289 =  ( n23 ) ? ( in_stream_buff_1 ) : ( n288 ) ;
assign n290 =  ( n18 ) ? ( in_stream_buff_1 ) : ( n289 ) ;
assign n291 =  ( n9 ) ? ( in_stream_buff_1 ) : ( n290 ) ;
assign n292 =  ( n4 ) ? ( in_stream_buff_1 ) : ( n291 ) ;
assign n293 =  ( in_stream_full ) == ( 1'd1 )  ;
assign n294 =  ( n293 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n295 =  ( n33 ) ? ( 1'd0 ) : ( in_stream_empty ) ;
assign n296 =  ( n28 ) ? ( n294 ) : ( n295 ) ;
assign n297 =  ( n23 ) ? ( in_stream_empty ) : ( n296 ) ;
assign n298 =  ( n18 ) ? ( in_stream_empty ) : ( n297 ) ;
assign n299 =  ( n9 ) ? ( in_stream_empty ) : ( n298 ) ;
assign n300 =  ( n4 ) ? ( in_stream_empty ) : ( n299 ) ;
assign n301 =  ( in_stream_empty ) == ( 1'd1 )  ;
assign n302 =  ( n301 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n303 =  ( n33 ) ? ( n302 ) : ( in_stream_full ) ;
assign n304 =  ( n28 ) ? ( 1'd0 ) : ( n303 ) ;
assign n305 =  ( n23 ) ? ( in_stream_full ) : ( n304 ) ;
assign n306 =  ( n18 ) ? ( in_stream_full ) : ( n305 ) ;
assign n307 =  ( n9 ) ? ( in_stream_full ) : ( n306 ) ;
assign n308 =  ( n4 ) ? ( in_stream_full ) : ( n307 ) ;
assign n309 =  ( n293 ) ? ( in_stream_buff_1 ) : ( in_stream_buff_0 ) ;
assign n310 =  ( LB2D_proc_w ) == ( 64'd0 )  ;
assign n311 =  (  LB2D_proc_7 [ LB2D_proc_x ] )  ;
assign n312 =  ( LB2D_proc_w ) == ( 64'd1 )  ;
assign n313 =  (  LB2D_proc_0 [ LB2D_proc_x ] )  ;
assign n314 =  ( LB2D_proc_w ) == ( 64'd2 )  ;
assign n315 =  (  LB2D_proc_1 [ LB2D_proc_x ] )  ;
assign n316 =  ( LB2D_proc_w ) == ( 64'd3 )  ;
assign n317 =  (  LB2D_proc_2 [ LB2D_proc_x ] )  ;
assign n318 =  ( LB2D_proc_w ) == ( 64'd4 )  ;
assign n319 =  (  LB2D_proc_3 [ LB2D_proc_x ] )  ;
assign n320 =  ( LB2D_proc_w ) == ( 64'd5 )  ;
assign n321 =  (  LB2D_proc_4 [ LB2D_proc_x ] )  ;
assign n322 =  ( LB2D_proc_w ) == ( 64'd6 )  ;
assign n323 =  (  LB2D_proc_5 [ LB2D_proc_x ] )  ;
assign n324 =  (  LB2D_proc_6 [ LB2D_proc_x ] )  ;
assign n325 =  ( n322 ) ? ( n323 ) : ( n324 ) ;
assign n326 =  ( n320 ) ? ( n321 ) : ( n325 ) ;
assign n327 =  ( n318 ) ? ( n319 ) : ( n326 ) ;
assign n328 =  ( n316 ) ? ( n317 ) : ( n327 ) ;
assign n329 =  ( n314 ) ? ( n315 ) : ( n328 ) ;
assign n330 =  ( n312 ) ? ( n313 ) : ( n329 ) ;
assign n331 =  ( n310 ) ? ( n311 ) : ( n330 ) ;
assign n332 =  ( n322 ) ? ( n321 ) : ( n323 ) ;
assign n333 =  ( n320 ) ? ( n319 ) : ( n332 ) ;
assign n334 =  ( n318 ) ? ( n317 ) : ( n333 ) ;
assign n335 =  ( n316 ) ? ( n315 ) : ( n334 ) ;
assign n336 =  ( n314 ) ? ( n313 ) : ( n335 ) ;
assign n337 =  ( n312 ) ? ( n311 ) : ( n336 ) ;
assign n338 =  ( n310 ) ? ( n324 ) : ( n337 ) ;
assign n339 =  ( n322 ) ? ( n319 ) : ( n321 ) ;
assign n340 =  ( n320 ) ? ( n317 ) : ( n339 ) ;
assign n341 =  ( n318 ) ? ( n315 ) : ( n340 ) ;
assign n342 =  ( n316 ) ? ( n313 ) : ( n341 ) ;
assign n343 =  ( n314 ) ? ( n311 ) : ( n342 ) ;
assign n344 =  ( n312 ) ? ( n324 ) : ( n343 ) ;
assign n345 =  ( n310 ) ? ( n323 ) : ( n344 ) ;
assign n346 =  ( n322 ) ? ( n317 ) : ( n319 ) ;
assign n347 =  ( n320 ) ? ( n315 ) : ( n346 ) ;
assign n348 =  ( n318 ) ? ( n313 ) : ( n347 ) ;
assign n349 =  ( n316 ) ? ( n311 ) : ( n348 ) ;
assign n350 =  ( n314 ) ? ( n324 ) : ( n349 ) ;
assign n351 =  ( n312 ) ? ( n323 ) : ( n350 ) ;
assign n352 =  ( n310 ) ? ( n321 ) : ( n351 ) ;
assign n353 =  ( n322 ) ? ( n315 ) : ( n317 ) ;
assign n354 =  ( n320 ) ? ( n313 ) : ( n353 ) ;
assign n355 =  ( n318 ) ? ( n311 ) : ( n354 ) ;
assign n356 =  ( n316 ) ? ( n324 ) : ( n355 ) ;
assign n357 =  ( n314 ) ? ( n323 ) : ( n356 ) ;
assign n358 =  ( n312 ) ? ( n321 ) : ( n357 ) ;
assign n359 =  ( n310 ) ? ( n319 ) : ( n358 ) ;
assign n360 =  ( n322 ) ? ( n313 ) : ( n315 ) ;
assign n361 =  ( n320 ) ? ( n311 ) : ( n360 ) ;
assign n362 =  ( n318 ) ? ( n324 ) : ( n361 ) ;
assign n363 =  ( n316 ) ? ( n323 ) : ( n362 ) ;
assign n364 =  ( n314 ) ? ( n321 ) : ( n363 ) ;
assign n365 =  ( n312 ) ? ( n319 ) : ( n364 ) ;
assign n366 =  ( n310 ) ? ( n317 ) : ( n365 ) ;
assign n367 =  ( n322 ) ? ( n311 ) : ( n313 ) ;
assign n368 =  ( n320 ) ? ( n324 ) : ( n367 ) ;
assign n369 =  ( n318 ) ? ( n323 ) : ( n368 ) ;
assign n370 =  ( n316 ) ? ( n321 ) : ( n369 ) ;
assign n371 =  ( n314 ) ? ( n319 ) : ( n370 ) ;
assign n372 =  ( n312 ) ? ( n317 ) : ( n371 ) ;
assign n373 =  ( n310 ) ? ( n315 ) : ( n372 ) ;
assign n374 =  ( n322 ) ? ( n324 ) : ( n311 ) ;
assign n375 =  ( n320 ) ? ( n323 ) : ( n374 ) ;
assign n376 =  ( n318 ) ? ( n321 ) : ( n375 ) ;
assign n377 =  ( n316 ) ? ( n319 ) : ( n376 ) ;
assign n378 =  ( n314 ) ? ( n317 ) : ( n377 ) ;
assign n379 =  ( n312 ) ? ( n315 ) : ( n378 ) ;
assign n380 =  ( n310 ) ? ( n313 ) : ( n379 ) ;
assign n381 =  { ( n373 ) , ( n380 ) }  ;
assign n382 =  { ( n366 ) , ( n381 ) }  ;
assign n383 =  { ( n359 ) , ( n382 ) }  ;
assign n384 =  { ( n352 ) , ( n383 ) }  ;
assign n385 =  { ( n345 ) , ( n384 ) }  ;
assign n386 =  { ( n338 ) , ( n385 ) }  ;
assign n387 =  { ( n331 ) , ( n386 ) }  ;
assign n388 =  { ( n309 ) , ( n387 ) }  ;
assign n389 =  ( n26 ) ? ( slice_stream_buff_0 ) : ( n388 ) ;
assign n390 =  ( n33 ) ? ( slice_stream_buff_0 ) : ( slice_stream_buff_0 ) ;
assign n391 =  ( n28 ) ? ( n389 ) : ( n390 ) ;
assign n392 =  ( n23 ) ? ( slice_stream_buff_0 ) : ( n391 ) ;
assign n393 =  ( n18 ) ? ( slice_stream_buff_0 ) : ( n392 ) ;
assign n394 =  ( n9 ) ? ( slice_stream_buff_0 ) : ( n393 ) ;
assign n395 =  ( n4 ) ? ( slice_stream_buff_0 ) : ( n394 ) ;
assign n396 =  ( n26 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n397 =  ( n33 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_1 ) ;
assign n398 =  ( n28 ) ? ( n396 ) : ( n397 ) ;
assign n399 =  ( n23 ) ? ( slice_stream_buff_1 ) : ( n398 ) ;
assign n400 =  ( n18 ) ? ( slice_stream_buff_1 ) : ( n399 ) ;
assign n401 =  ( n9 ) ? ( slice_stream_buff_1 ) : ( n400 ) ;
assign n402 =  ( n4 ) ? ( slice_stream_buff_1 ) : ( n401 ) ;
assign n403 =  ( n76 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n404 =  ( n26 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n405 =  ( n33 ) ? ( slice_stream_empty ) : ( slice_stream_empty ) ;
assign n406 =  ( n28 ) ? ( n404 ) : ( n405 ) ;
assign n407 =  ( n23 ) ? ( n403 ) : ( n406 ) ;
assign n408 =  ( n18 ) ? ( slice_stream_empty ) : ( n407 ) ;
assign n409 =  ( n9 ) ? ( slice_stream_empty ) : ( n408 ) ;
assign n410 =  ( n4 ) ? ( slice_stream_empty ) : ( n409 ) ;
assign n411 =  ( slice_stream_empty ) == ( 1'd1 )  ;
assign n412 =  ( n411 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n413 =  ( n26 ) ? ( 1'd0 ) : ( n412 ) ;
assign n414 =  ( n33 ) ? ( slice_stream_full ) : ( slice_stream_full ) ;
assign n415 =  ( n28 ) ? ( n413 ) : ( n414 ) ;
assign n416 =  ( n23 ) ? ( 1'd0 ) : ( n415 ) ;
assign n417 =  ( n18 ) ? ( slice_stream_full ) : ( n416 ) ;
assign n418 =  ( n9 ) ? ( slice_stream_full ) : ( n417 ) ;
assign n419 =  ( n4 ) ? ( slice_stream_full ) : ( n418 ) ;
assign n420 =  ( LB2D_shift_x ) >= ( 9'd8 )  ;
assign n421 = n77[71:64] ;
assign n422 = LB2D_shift_0[71:64] ;
assign n423 = LB2D_shift_1[71:64] ;
assign n424 = LB2D_shift_2[71:64] ;
assign n425 = LB2D_shift_3[71:64] ;
assign n426 = LB2D_shift_4[71:64] ;
assign n427 = LB2D_shift_5[71:64] ;
assign n428 = LB2D_shift_6[71:64] ;
assign n429 = LB2D_shift_7[71:64] ;
assign n430 =  { ( n428 ) , ( n429 ) }  ;
assign n431 =  { ( n427 ) , ( n430 ) }  ;
assign n432 =  { ( n426 ) , ( n431 ) }  ;
assign n433 =  { ( n425 ) , ( n432 ) }  ;
assign n434 =  { ( n424 ) , ( n433 ) }  ;
assign n435 =  { ( n423 ) , ( n434 ) }  ;
assign n436 =  { ( n422 ) , ( n435 ) }  ;
assign n437 =  { ( n421 ) , ( n436 ) }  ;
assign n438 = n77[63:56] ;
assign n439 = LB2D_shift_0[63:56] ;
assign n440 = LB2D_shift_1[63:56] ;
assign n441 = LB2D_shift_2[63:56] ;
assign n442 = LB2D_shift_3[63:56] ;
assign n443 = LB2D_shift_4[63:56] ;
assign n444 = LB2D_shift_5[63:56] ;
assign n445 = LB2D_shift_6[63:56] ;
assign n446 = LB2D_shift_7[63:56] ;
assign n447 =  { ( n445 ) , ( n446 ) }  ;
assign n448 =  { ( n444 ) , ( n447 ) }  ;
assign n449 =  { ( n443 ) , ( n448 ) }  ;
assign n450 =  { ( n442 ) , ( n449 ) }  ;
assign n451 =  { ( n441 ) , ( n450 ) }  ;
assign n452 =  { ( n440 ) , ( n451 ) }  ;
assign n453 =  { ( n439 ) , ( n452 ) }  ;
assign n454 =  { ( n438 ) , ( n453 ) }  ;
assign n455 = n77[55:48] ;
assign n456 = LB2D_shift_0[55:48] ;
assign n457 = LB2D_shift_1[55:48] ;
assign n458 = LB2D_shift_2[55:48] ;
assign n459 = LB2D_shift_3[55:48] ;
assign n460 = LB2D_shift_4[55:48] ;
assign n461 = LB2D_shift_5[55:48] ;
assign n462 = LB2D_shift_6[55:48] ;
assign n463 = LB2D_shift_7[55:48] ;
assign n464 =  { ( n462 ) , ( n463 ) }  ;
assign n465 =  { ( n461 ) , ( n464 ) }  ;
assign n466 =  { ( n460 ) , ( n465 ) }  ;
assign n467 =  { ( n459 ) , ( n466 ) }  ;
assign n468 =  { ( n458 ) , ( n467 ) }  ;
assign n469 =  { ( n457 ) , ( n468 ) }  ;
assign n470 =  { ( n456 ) , ( n469 ) }  ;
assign n471 =  { ( n455 ) , ( n470 ) }  ;
assign n472 = n77[47:40] ;
assign n473 = LB2D_shift_0[47:40] ;
assign n474 = LB2D_shift_1[47:40] ;
assign n475 = LB2D_shift_2[47:40] ;
assign n476 = LB2D_shift_3[47:40] ;
assign n477 = LB2D_shift_4[47:40] ;
assign n478 = LB2D_shift_5[47:40] ;
assign n479 = LB2D_shift_6[47:40] ;
assign n480 = LB2D_shift_7[47:40] ;
assign n481 =  { ( n479 ) , ( n480 ) }  ;
assign n482 =  { ( n478 ) , ( n481 ) }  ;
assign n483 =  { ( n477 ) , ( n482 ) }  ;
assign n484 =  { ( n476 ) , ( n483 ) }  ;
assign n485 =  { ( n475 ) , ( n484 ) }  ;
assign n486 =  { ( n474 ) , ( n485 ) }  ;
assign n487 =  { ( n473 ) , ( n486 ) }  ;
assign n488 =  { ( n472 ) , ( n487 ) }  ;
assign n489 = n77[39:32] ;
assign n490 = LB2D_shift_0[39:32] ;
assign n491 = LB2D_shift_1[39:32] ;
assign n492 = LB2D_shift_2[39:32] ;
assign n493 = LB2D_shift_3[39:32] ;
assign n494 = LB2D_shift_4[39:32] ;
assign n495 = LB2D_shift_5[39:32] ;
assign n496 = LB2D_shift_6[39:32] ;
assign n497 = LB2D_shift_7[39:32] ;
assign n498 =  { ( n496 ) , ( n497 ) }  ;
assign n499 =  { ( n495 ) , ( n498 ) }  ;
assign n500 =  { ( n494 ) , ( n499 ) }  ;
assign n501 =  { ( n493 ) , ( n500 ) }  ;
assign n502 =  { ( n492 ) , ( n501 ) }  ;
assign n503 =  { ( n491 ) , ( n502 ) }  ;
assign n504 =  { ( n490 ) , ( n503 ) }  ;
assign n505 =  { ( n489 ) , ( n504 ) }  ;
assign n506 = n77[31:24] ;
assign n507 = LB2D_shift_0[31:24] ;
assign n508 = LB2D_shift_1[31:24] ;
assign n509 = LB2D_shift_2[31:24] ;
assign n510 = LB2D_shift_3[31:24] ;
assign n511 = LB2D_shift_4[31:24] ;
assign n512 = LB2D_shift_5[31:24] ;
assign n513 = LB2D_shift_6[31:24] ;
assign n514 = LB2D_shift_7[31:24] ;
assign n515 =  { ( n513 ) , ( n514 ) }  ;
assign n516 =  { ( n512 ) , ( n515 ) }  ;
assign n517 =  { ( n511 ) , ( n516 ) }  ;
assign n518 =  { ( n510 ) , ( n517 ) }  ;
assign n519 =  { ( n509 ) , ( n518 ) }  ;
assign n520 =  { ( n508 ) , ( n519 ) }  ;
assign n521 =  { ( n507 ) , ( n520 ) }  ;
assign n522 =  { ( n506 ) , ( n521 ) }  ;
assign n523 = n77[23:16] ;
assign n524 = LB2D_shift_0[23:16] ;
assign n525 = LB2D_shift_1[23:16] ;
assign n526 = LB2D_shift_2[23:16] ;
assign n527 = LB2D_shift_3[23:16] ;
assign n528 = LB2D_shift_4[23:16] ;
assign n529 = LB2D_shift_5[23:16] ;
assign n530 = LB2D_shift_6[23:16] ;
assign n531 = LB2D_shift_7[23:16] ;
assign n532 =  { ( n530 ) , ( n531 ) }  ;
assign n533 =  { ( n529 ) , ( n532 ) }  ;
assign n534 =  { ( n528 ) , ( n533 ) }  ;
assign n535 =  { ( n527 ) , ( n534 ) }  ;
assign n536 =  { ( n526 ) , ( n535 ) }  ;
assign n537 =  { ( n525 ) , ( n536 ) }  ;
assign n538 =  { ( n524 ) , ( n537 ) }  ;
assign n539 =  { ( n523 ) , ( n538 ) }  ;
assign n540 = n77[15:8] ;
assign n541 = LB2D_shift_0[15:8] ;
assign n542 = LB2D_shift_1[15:8] ;
assign n543 = LB2D_shift_2[15:8] ;
assign n544 = LB2D_shift_3[15:8] ;
assign n545 = LB2D_shift_4[15:8] ;
assign n546 = LB2D_shift_5[15:8] ;
assign n547 = LB2D_shift_6[15:8] ;
assign n548 = LB2D_shift_7[15:8] ;
assign n549 =  { ( n547 ) , ( n548 ) }  ;
assign n550 =  { ( n546 ) , ( n549 ) }  ;
assign n551 =  { ( n545 ) , ( n550 ) }  ;
assign n552 =  { ( n544 ) , ( n551 ) }  ;
assign n553 =  { ( n543 ) , ( n552 ) }  ;
assign n554 =  { ( n542 ) , ( n553 ) }  ;
assign n555 =  { ( n541 ) , ( n554 ) }  ;
assign n556 =  { ( n540 ) , ( n555 ) }  ;
assign n557 = n77[7:0] ;
assign n558 = LB2D_shift_0[7:0] ;
assign n559 = LB2D_shift_1[7:0] ;
assign n560 = LB2D_shift_2[7:0] ;
assign n561 = LB2D_shift_3[7:0] ;
assign n562 = LB2D_shift_4[7:0] ;
assign n563 = LB2D_shift_5[7:0] ;
assign n564 = LB2D_shift_6[7:0] ;
assign n565 = LB2D_shift_7[7:0] ;
assign n566 =  { ( n564 ) , ( n565 ) }  ;
assign n567 =  { ( n563 ) , ( n566 ) }  ;
assign n568 =  { ( n562 ) , ( n567 ) }  ;
assign n569 =  { ( n561 ) , ( n568 ) }  ;
assign n570 =  { ( n560 ) , ( n569 ) }  ;
assign n571 =  { ( n559 ) , ( n570 ) }  ;
assign n572 =  { ( n558 ) , ( n571 ) }  ;
assign n573 =  { ( n557 ) , ( n572 ) }  ;
assign n574 =  { ( n556 ) , ( n573 ) }  ;
assign n575 =  { ( n539 ) , ( n574 ) }  ;
assign n576 =  { ( n522 ) , ( n575 ) }  ;
assign n577 =  { ( n505 ) , ( n576 ) }  ;
assign n578 =  { ( n488 ) , ( n577 ) }  ;
assign n579 =  { ( n471 ) , ( n578 ) }  ;
assign n580 =  { ( n454 ) , ( n579 ) }  ;
assign n581 =  { ( n437 ) , ( n580 ) }  ;
assign n582 =  ( n420 ) ? ( n581 ) : ( stencil_stream_buff_0 ) ;
assign n583 =  ( n33 ) ? ( stencil_stream_buff_0 ) : ( stencil_stream_buff_0 ) ;
assign n584 =  ( n28 ) ? ( stencil_stream_buff_0 ) : ( n583 ) ;
assign n585 =  ( n23 ) ? ( n582 ) : ( n584 ) ;
assign n586 =  ( n18 ) ? ( stencil_stream_buff_0 ) : ( n585 ) ;
assign n587 =  ( n9 ) ? ( stencil_stream_buff_0 ) : ( n586 ) ;
assign n588 =  ( n4 ) ? ( stencil_stream_buff_0 ) : ( n587 ) ;
assign n589 =  ( n33 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_1 ) ;
assign n590 =  ( n28 ) ? ( stencil_stream_buff_1 ) : ( n589 ) ;
assign n591 =  ( n23 ) ? ( stencil_stream_buff_0 ) : ( n590 ) ;
assign n592 =  ( n18 ) ? ( stencil_stream_buff_1 ) : ( n591 ) ;
assign n593 =  ( n9 ) ? ( stencil_stream_buff_1 ) : ( n592 ) ;
assign n594 =  ( n4 ) ? ( stencil_stream_buff_1 ) : ( n593 ) ;
assign n595 =  ( n145 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n596 =  ( n21 ) ? ( stencil_stream_empty ) : ( 1'd0 ) ;
assign n597 =  ( n33 ) ? ( stencil_stream_empty ) : ( stencil_stream_empty ) ;
assign n598 =  ( n28 ) ? ( stencil_stream_empty ) : ( n597 ) ;
assign n599 =  ( n23 ) ? ( n596 ) : ( n598 ) ;
assign n600 =  ( n18 ) ? ( n595 ) : ( n599 ) ;
assign n601 =  ( n9 ) ? ( stencil_stream_empty ) : ( n600 ) ;
assign n602 =  ( n4 ) ? ( stencil_stream_empty ) : ( n601 ) ;
assign n603 =  ( n14 ) ? ( 1'd0 ) : ( 1'd0 ) ;
assign n604 =  ( stencil_stream_empty ) == ( 1'd1 )  ;
assign n605 =  ( n604 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n606 =  ( n21 ) ? ( stencil_stream_full ) : ( n605 ) ;
assign n607 =  ( n33 ) ? ( stencil_stream_full ) : ( stencil_stream_full ) ;
assign n608 =  ( n28 ) ? ( stencil_stream_full ) : ( n607 ) ;
assign n609 =  ( n23 ) ? ( n606 ) : ( n608 ) ;
assign n610 =  ( n18 ) ? ( n603 ) : ( n609 ) ;
assign n611 =  ( n9 ) ? ( stencil_stream_full ) : ( n610 ) ;
assign n612 =  ( n4 ) ? ( stencil_stream_full ) : ( n611 ) ;
assign n613 = ~ ( n4 ) ;
assign n614 = ~ ( n9 ) ;
assign n615 =  ( n613 ) & ( n614 )  ;
assign n616 = ~ ( n18 ) ;
assign n617 =  ( n615 ) & ( n616 )  ;
assign n618 = ~ ( n23 ) ;
assign n619 =  ( n617 ) & ( n618 )  ;
assign n620 = ~ ( n28 ) ;
assign n621 =  ( n619 ) & ( n620 )  ;
assign n622 = ~ ( n33 ) ;
assign n623 =  ( n621 ) & ( n622 )  ;
assign n624 =  ( n621 ) & ( n33 )  ;
assign n625 =  ( n619 ) & ( n28 )  ;
assign n626 = ~ ( n310 ) ;
assign n627 =  ( n625 ) & ( n626 )  ;
assign n628 =  ( n625 ) & ( n310 )  ;
assign n629 =  ( n617 ) & ( n23 )  ;
assign n630 =  ( n615 ) & ( n18 )  ;
assign n631 =  ( n613 ) & ( n9 )  ;
assign LB2D_proc_0_addr0 = n628 ? (LB2D_proc_x) : (0);
assign LB2D_proc_0_data0 = n628 ? (n309) : (LB2D_proc_0[0]);
assign n632 = ~ ( n312 ) ;
assign n633 =  ( n625 ) & ( n632 )  ;
assign n634 =  ( n625 ) & ( n312 )  ;
assign LB2D_proc_1_addr0 = n634 ? (LB2D_proc_x) : (0);
assign LB2D_proc_1_data0 = n634 ? (n309) : (LB2D_proc_1[0]);
assign n635 = ~ ( n314 ) ;
assign n636 =  ( n625 ) & ( n635 )  ;
assign n637 =  ( n625 ) & ( n314 )  ;
assign LB2D_proc_2_addr0 = n637 ? (LB2D_proc_x) : (0);
assign LB2D_proc_2_data0 = n637 ? (n309) : (LB2D_proc_2[0]);
assign n638 = ~ ( n316 ) ;
assign n639 =  ( n625 ) & ( n638 )  ;
assign n640 =  ( n625 ) & ( n316 )  ;
assign LB2D_proc_3_addr0 = n640 ? (LB2D_proc_x) : (0);
assign LB2D_proc_3_data0 = n640 ? (n309) : (LB2D_proc_3[0]);
assign n641 = ~ ( n318 ) ;
assign n642 =  ( n625 ) & ( n641 )  ;
assign n643 =  ( n625 ) & ( n318 )  ;
assign LB2D_proc_4_addr0 = n643 ? (LB2D_proc_x) : (0);
assign LB2D_proc_4_data0 = n643 ? (n309) : (LB2D_proc_4[0]);
assign n644 = ~ ( n320 ) ;
assign n645 =  ( n625 ) & ( n644 )  ;
assign n646 =  ( n625 ) & ( n320 )  ;
assign LB2D_proc_5_addr0 = n646 ? (LB2D_proc_x) : (0);
assign LB2D_proc_5_data0 = n646 ? (n309) : (LB2D_proc_5[0]);
assign n647 = ~ ( n322 ) ;
assign n648 =  ( n625 ) & ( n647 )  ;
assign n649 =  ( n625 ) & ( n322 )  ;
assign LB2D_proc_6_addr0 = n649 ? (LB2D_proc_x) : (0);
assign LB2D_proc_6_data0 = n649 ? (n309) : (LB2D_proc_6[0]);
assign n650 =  ( LB2D_proc_w ) == ( 64'd7 )  ;
assign n651 = ~ ( n650 ) ;
assign n652 =  ( n625 ) & ( n651 )  ;
assign n653 =  ( n625 ) & ( n650 )  ;
assign LB2D_proc_7_addr0 = n653 ? (LB2D_proc_x) : (0);
assign LB2D_proc_7_data0 = n653 ? (n309) : (LB2D_proc_7[0]);
/*
function [7:0] gb_fun ;
input [647:0] arg0;
    begin
//TODO: Add the specific function HERE.    end
endfunction
*/

always @(posedge clk) begin
   if(rst) begin
       LB1D_buff <= LB1D_buff;
       LB1D_p_cnt <= LB1D_p_cnt;
       LB2D_proc_w <= LB2D_proc_w;
       LB2D_proc_x <= LB2D_proc_x;
       LB2D_proc_y <= LB2D_proc_y;
       LB2D_shift_0 <= LB2D_shift_0;
       LB2D_shift_1 <= LB2D_shift_1;
       LB2D_shift_2 <= LB2D_shift_2;
       LB2D_shift_3 <= LB2D_shift_3;
       LB2D_shift_4 <= LB2D_shift_4;
       LB2D_shift_5 <= LB2D_shift_5;
       LB2D_shift_6 <= LB2D_shift_6;
       LB2D_shift_7 <= LB2D_shift_7;
       LB2D_shift_x <= LB2D_shift_x;
       LB2D_shift_y <= LB2D_shift_y;
       arg_0_TDATA <= arg_0_TDATA;
       arg_0_TVALID <= arg_0_TVALID;
       arg_1_TREADY <= arg_1_TREADY;
       gb_exit_it_1 <= gb_exit_it_1;
       gb_exit_it_2 <= gb_exit_it_2;
       gb_exit_it_3 <= gb_exit_it_3;
       gb_exit_it_4 <= gb_exit_it_4;
       gb_exit_it_5 <= gb_exit_it_5;
       gb_exit_it_6 <= gb_exit_it_6;
       gb_exit_it_7 <= gb_exit_it_7;
       gb_exit_it_8 <= gb_exit_it_8;
       gb_p_cnt <= gb_p_cnt;
       gb_pp_it_1 <= gb_pp_it_1;
       gb_pp_it_2 <= gb_pp_it_2;
       gb_pp_it_3 <= gb_pp_it_3;
       gb_pp_it_4 <= gb_pp_it_4;
       gb_pp_it_5 <= gb_pp_it_5;
       gb_pp_it_6 <= gb_pp_it_6;
       gb_pp_it_7 <= gb_pp_it_7;
       gb_pp_it_8 <= gb_pp_it_8;
       gb_pp_it_9 <= gb_pp_it_9;
       in_stream_buff_0 <= in_stream_buff_0;
       in_stream_buff_1 <= in_stream_buff_1;
       in_stream_empty <= in_stream_empty;
       in_stream_full <= in_stream_full;
       slice_stream_buff_0 <= slice_stream_buff_0;
       slice_stream_buff_1 <= slice_stream_buff_1;
       slice_stream_empty <= slice_stream_empty;
       slice_stream_full <= slice_stream_full;
       stencil_stream_buff_0 <= stencil_stream_buff_0;
       stencil_stream_buff_1 <= stencil_stream_buff_1;
       stencil_stream_empty <= stencil_stream_empty;
       stencil_stream_full <= stencil_stream_full;
   end
   else if(step) begin
       LB1D_buff <= n39;
       LB1D_p_cnt <= n46;
       LB2D_proc_w <= n57;
       LB2D_proc_x <= n65;
       LB2D_proc_y <= n75;
       LB2D_shift_0 <= n83;
       LB2D_shift_1 <= n89;
       LB2D_shift_2 <= n95;
       LB2D_shift_3 <= n101;
       LB2D_shift_4 <= n107;
       LB2D_shift_5 <= n113;
       LB2D_shift_6 <= n119;
       LB2D_shift_7 <= n125;
       LB2D_shift_x <= n134;
       LB2D_shift_y <= n144;
       arg_0_TDATA <= n153;
       arg_0_TVALID <= n161;
       arg_1_TREADY <= n167;
       gb_exit_it_1 <= n176;
       gb_exit_it_2 <= n182;
       gb_exit_it_3 <= n188;
       gb_exit_it_4 <= n194;
       gb_exit_it_5 <= n200;
       gb_exit_it_6 <= n206;
       gb_exit_it_7 <= n212;
       gb_exit_it_8 <= n218;
       gb_p_cnt <= n226;
       gb_pp_it_1 <= n232;
       gb_pp_it_2 <= n238;
       gb_pp_it_3 <= n244;
       gb_pp_it_4 <= n250;
       gb_pp_it_5 <= n256;
       gb_pp_it_6 <= n262;
       gb_pp_it_7 <= n268;
       gb_pp_it_8 <= n274;
       gb_pp_it_9 <= n280;
       in_stream_buff_0 <= n286;
       in_stream_buff_1 <= n292;
       in_stream_empty <= n300;
       in_stream_full <= n308;
       slice_stream_buff_0 <= n395;
       slice_stream_buff_1 <= n402;
       slice_stream_empty <= n410;
       slice_stream_full <= n419;
       stencil_stream_buff_0 <= n588;
       stencil_stream_buff_1 <= n594;
       stencil_stream_empty <= n602;
       stencil_stream_full <= n612;
       LB2D_proc_0 [ LB2D_proc_0_addr0 ] <= LB2D_proc_0_data0;
       LB2D_proc_1 [ LB2D_proc_1_addr0 ] <= LB2D_proc_1_data0;
       LB2D_proc_2 [ LB2D_proc_2_addr0 ] <= LB2D_proc_2_data0;
       LB2D_proc_3 [ LB2D_proc_3_addr0 ] <= LB2D_proc_3_data0;
       LB2D_proc_4 [ LB2D_proc_4_addr0 ] <= LB2D_proc_4_data0;
       LB2D_proc_5 [ LB2D_proc_5_addr0 ] <= LB2D_proc_5_data0;
       LB2D_proc_6 [ LB2D_proc_6_addr0 ] <= LB2D_proc_6_data0;
       LB2D_proc_7 [ LB2D_proc_7_addr0 ] <= LB2D_proc_7_data0;
   end
end
endmodule
