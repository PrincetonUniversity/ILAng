module GB(
arg_0_TREADY,
arg_1_TDATA,
arg_1_TVALID,
LB1D_buff,
LB1D_in,
LB1D_it_1,
LB1D_p_cnt,
LB2D_proc_w,
LB2D_proc_x,
LB2D_proc_y,
LB2D_shift_0,
LB2D_shift_1,
LB2D_shift_2,
LB2D_shift_3,
LB2D_shift_4,
LB2D_shift_5,
LB2D_shift_6,
LB2D_shift_7,
LB2D_shift_x,
LB2D_shift_y,
arg_0_TDATA,
arg_0_TVALID,
arg_1_TREADY,
gb_exit_it_1,
gb_exit_it_2,
gb_exit_it_3,
gb_exit_it_4,
gb_exit_it_5,
gb_exit_it_6,
gb_exit_it_7,
gb_exit_it_8,
gb_p_cnt,
gb_pp_it_1,
gb_pp_it_2,
gb_pp_it_3,
gb_pp_it_4,
gb_pp_it_5,
gb_pp_it_6,
gb_pp_it_7,
gb_pp_it_8,
gb_pp_it_9,
in_stream_buff_0,
in_stream_buff_1,
in_stream_empty,
in_stream_full,
slice_stream_buff_0,
slice_stream_buff_1,
slice_stream_empty,
slice_stream_full,
stencil_stream_buff_0,
stencil_stream_buff_1,
stencil_stream_empty,
stencil_stream_full,
clk,rst,
step
);
input            arg_0_TREADY;
input      [7:0] arg_1_TDATA;
input            arg_1_TVALID;
input clk;
input rst;
input step;
output      [7:0] LB1D_buff;
output      [7:0] LB1D_in;
output            LB1D_it_1;
output     [18:0] LB1D_p_cnt;
output     [63:0] LB2D_proc_w;
output      [8:0] LB2D_proc_x;
output      [9:0] LB2D_proc_y;
output     [71:0] LB2D_shift_0;
output     [71:0] LB2D_shift_1;
output     [71:0] LB2D_shift_2;
output     [71:0] LB2D_shift_3;
output     [71:0] LB2D_shift_4;
output     [71:0] LB2D_shift_5;
output     [71:0] LB2D_shift_6;
output     [71:0] LB2D_shift_7;
output      [8:0] LB2D_shift_x;
output      [9:0] LB2D_shift_y;
output      [7:0] arg_0_TDATA;
output            arg_0_TVALID;
output            arg_1_TREADY;
output            gb_exit_it_1;
output            gb_exit_it_2;
output            gb_exit_it_3;
output            gb_exit_it_4;
output            gb_exit_it_5;
output            gb_exit_it_6;
output            gb_exit_it_7;
output            gb_exit_it_8;
output     [18:0] gb_p_cnt;
output            gb_pp_it_1;
output            gb_pp_it_2;
output            gb_pp_it_3;
output            gb_pp_it_4;
output            gb_pp_it_5;
output            gb_pp_it_6;
output            gb_pp_it_7;
output            gb_pp_it_8;
output            gb_pp_it_9;
output      [7:0] in_stream_buff_0;
output      [7:0] in_stream_buff_1;
output            in_stream_empty;
output            in_stream_full;
output     [71:0] slice_stream_buff_0;
output     [71:0] slice_stream_buff_1;
output            slice_stream_empty;
output            slice_stream_full;
output    [647:0] stencil_stream_buff_0;
output    [647:0] stencil_stream_buff_1;
output            stencil_stream_empty;
output            stencil_stream_full;
reg      [7:0] LB1D_buff;
reg      [7:0] LB1D_in;
reg            LB1D_it_1;
reg     [18:0] LB1D_p_cnt;
reg     [63:0] LB2D_proc_w;
reg      [8:0] LB2D_proc_x;
reg      [9:0] LB2D_proc_y;
reg     [71:0] LB2D_shift_0;
reg     [71:0] LB2D_shift_1;
reg     [71:0] LB2D_shift_2;
reg     [71:0] LB2D_shift_3;
reg     [71:0] LB2D_shift_4;
reg     [71:0] LB2D_shift_5;
reg     [71:0] LB2D_shift_6;
reg     [71:0] LB2D_shift_7;
reg      [8:0] LB2D_shift_x;
reg      [9:0] LB2D_shift_y;
reg      [7:0] arg_0_TDATA;
reg            arg_0_TVALID;
reg            arg_1_TREADY;
reg            gb_exit_it_1;
reg            gb_exit_it_2;
reg            gb_exit_it_3;
reg            gb_exit_it_4;
reg            gb_exit_it_5;
reg            gb_exit_it_6;
reg            gb_exit_it_7;
reg            gb_exit_it_8;
reg     [18:0] gb_p_cnt;
reg            gb_pp_it_1;
reg            gb_pp_it_2;
reg            gb_pp_it_3;
reg            gb_pp_it_4;
reg            gb_pp_it_5;
reg            gb_pp_it_6;
reg            gb_pp_it_7;
reg            gb_pp_it_8;
reg            gb_pp_it_9;
reg      [7:0] in_stream_buff_0;
reg      [7:0] in_stream_buff_1;
reg            in_stream_empty;
reg            in_stream_full;
reg     [71:0] slice_stream_buff_0;
reg     [71:0] slice_stream_buff_1;
reg            slice_stream_empty;
reg            slice_stream_full;
reg    [647:0] stencil_stream_buff_0;
reg    [647:0] stencil_stream_buff_1;
reg            stencil_stream_empty;
reg            stencil_stream_full;
wire            arg_0_TREADY;
wire      [7:0] arg_1_TDATA;
wire            arg_1_TVALID;
wire            n0;
wire            n1;
wire            n2;
wire            n3;
wire            n4;
wire            n5;
wire            n6;
wire            n7;
wire            n8;
wire            n9;
wire            n10;
wire            n11;
wire            n12;
wire            n13;
wire            n14;
wire            n15;
wire            n16;
wire            n17;
wire            n18;
wire            n19;
wire            n20;
wire            n21;
wire            n22;
wire            n23;
wire            n24;
wire            n25;
wire            n26;
wire            n27;
wire            n28;
wire            n29;
wire            n30;
wire      [7:0] n31;
wire      [7:0] n32;
wire      [7:0] n33;
wire      [7:0] n34;
wire      [7:0] n35;
wire      [7:0] n36;
wire      [7:0] n37;
wire      [7:0] n38;
wire      [7:0] n39;
wire            n40;
wire            n41;
wire            n42;
wire            n43;
wire            n44;
wire            n45;
wire            n46;
wire            n47;
wire            n48;
wire            n49;
wire     [18:0] n50;
wire     [18:0] n51;
wire            n52;
wire     [18:0] n53;
wire     [18:0] n54;
wire     [18:0] n55;
wire     [18:0] n56;
wire     [18:0] n57;
wire     [18:0] n58;
wire     [18:0] n59;
wire     [18:0] n60;
wire            n61;
wire            n62;
wire     [63:0] n63;
wire     [63:0] n64;
wire     [63:0] n65;
wire     [63:0] n66;
wire     [63:0] n67;
wire     [63:0] n68;
wire     [63:0] n69;
wire     [63:0] n70;
wire     [63:0] n71;
wire            n72;
wire            n73;
wire            n74;
wire      [8:0] n75;
wire      [8:0] n76;
wire      [8:0] n77;
wire      [8:0] n78;
wire      [8:0] n79;
wire      [8:0] n80;
wire      [8:0] n81;
wire      [8:0] n82;
wire            n83;
wire      [9:0] n84;
wire      [9:0] n85;
wire      [9:0] n86;
wire      [9:0] n87;
wire      [9:0] n88;
wire      [9:0] n89;
wire      [9:0] n90;
wire            n91;
wire     [71:0] n92;
wire     [71:0] n93;
wire     [71:0] n94;
wire     [71:0] n95;
wire     [71:0] n96;
wire     [71:0] n97;
wire     [71:0] n98;
wire     [71:0] n99;
wire     [71:0] n100;
wire     [71:0] n101;
wire     [71:0] n102;
wire     [71:0] n103;
wire     [71:0] n104;
wire     [71:0] n105;
wire     [71:0] n106;
wire     [71:0] n107;
wire     [71:0] n108;
wire     [71:0] n109;
wire     [71:0] n110;
wire     [71:0] n111;
wire     [71:0] n112;
wire     [71:0] n113;
wire     [71:0] n114;
wire     [71:0] n115;
wire     [71:0] n116;
wire     [71:0] n117;
wire     [71:0] n118;
wire     [71:0] n119;
wire     [71:0] n120;
wire     [71:0] n121;
wire     [71:0] n122;
wire     [71:0] n123;
wire     [71:0] n124;
wire     [71:0] n125;
wire     [71:0] n126;
wire     [71:0] n127;
wire     [71:0] n128;
wire     [71:0] n129;
wire     [71:0] n130;
wire     [71:0] n131;
wire     [71:0] n132;
wire     [71:0] n133;
wire     [71:0] n134;
wire     [71:0] n135;
wire     [71:0] n136;
wire     [71:0] n137;
wire     [71:0] n138;
wire     [71:0] n139;
wire     [71:0] n140;
wire      [8:0] n141;
wire      [8:0] n142;
wire      [8:0] n143;
wire      [8:0] n144;
wire      [8:0] n145;
wire      [8:0] n146;
wire      [8:0] n147;
wire            n148;
wire            n149;
wire      [9:0] n150;
wire      [9:0] n151;
wire      [9:0] n152;
wire      [9:0] n153;
wire      [9:0] n154;
wire      [9:0] n155;
wire      [9:0] n156;
wire      [9:0] n157;
wire      [9:0] n158;
wire            n159;
wire    [647:0] n160;
wire      [7:0] n161;
wire      [7:0] n162;
wire      [7:0] n163;
wire      [7:0] n164;
wire      [7:0] n165;
wire      [7:0] n166;
wire      [7:0] n167;
wire            n168;
wire            n169;
wire            n170;
wire            n171;
wire            n172;
wire            n173;
wire            n174;
wire            n175;
wire            n176;
wire            n177;
wire            n178;
wire            n179;
wire            n180;
wire            n181;
wire            n182;
wire     [18:0] n183;
wire            n184;
wire            n185;
wire            n186;
wire            n187;
wire            n188;
wire            n189;
wire            n190;
wire            n191;
wire            n192;
wire            n193;
wire            n194;
wire            n195;
wire            n196;
wire            n197;
wire            n198;
wire            n199;
wire            n200;
wire            n201;
wire            n202;
wire            n203;
wire            n204;
wire            n205;
wire            n206;
wire            n207;
wire            n208;
wire            n209;
wire            n210;
wire            n211;
wire            n212;
wire            n213;
wire            n214;
wire            n215;
wire            n216;
wire            n217;
wire            n218;
wire            n219;
wire            n220;
wire            n221;
wire            n222;
wire            n223;
wire            n224;
wire            n225;
wire            n226;
wire            n227;
wire            n228;
wire            n229;
wire            n230;
wire            n231;
wire            n232;
wire            n233;
wire            n234;
wire     [18:0] n235;
wire     [18:0] n236;
wire     [18:0] n237;
wire     [18:0] n238;
wire     [18:0] n239;
wire     [18:0] n240;
wire     [18:0] n241;
wire            n242;
wire            n243;
wire            n244;
wire            n245;
wire            n246;
wire            n247;
wire            n248;
wire            n249;
wire            n250;
wire            n251;
wire            n252;
wire            n253;
wire            n254;
wire            n255;
wire            n256;
wire            n257;
wire            n258;
wire            n259;
wire            n260;
wire            n261;
wire            n262;
wire            n263;
wire            n264;
wire            n265;
wire            n266;
wire            n267;
wire            n268;
wire            n269;
wire            n270;
wire            n271;
wire            n272;
wire            n273;
wire            n274;
wire            n275;
wire            n276;
wire            n277;
wire            n278;
wire            n279;
wire            n280;
wire            n281;
wire            n282;
wire            n283;
wire            n284;
wire            n285;
wire            n286;
wire            n287;
wire            n288;
wire            n289;
wire            n290;
wire            n291;
wire            n292;
wire            n293;
wire            n294;
wire            n295;
wire      [7:0] n296;
wire      [7:0] n297;
wire      [7:0] n298;
wire      [7:0] n299;
wire      [7:0] n300;
wire      [7:0] n301;
wire      [7:0] n302;
wire      [7:0] n303;
wire      [7:0] n304;
wire      [7:0] n305;
wire      [7:0] n306;
wire      [7:0] n307;
wire            n308;
wire            n309;
wire            n310;
wire            n311;
wire            n312;
wire            n313;
wire            n314;
wire            n315;
wire            n316;
wire            n317;
wire            n318;
wire            n319;
wire            n320;
wire            n321;
wire            n322;
wire            n323;
wire      [7:0] n324;
wire            n325;
wire      [7:0] n326;
wire            n327;
wire      [7:0] n328;
wire            n329;
wire      [7:0] n330;
wire            n331;
wire      [7:0] n332;
wire            n333;
wire      [7:0] n334;
wire            n335;
wire      [7:0] n336;
wire            n337;
wire      [7:0] n338;
wire      [7:0] n339;
wire      [7:0] n340;
wire      [7:0] n341;
wire      [7:0] n342;
wire      [7:0] n343;
wire      [7:0] n344;
wire      [7:0] n345;
wire      [7:0] n346;
wire      [7:0] n347;
wire      [7:0] n348;
wire      [7:0] n349;
wire      [7:0] n350;
wire      [7:0] n351;
wire      [7:0] n352;
wire      [7:0] n353;
wire      [7:0] n354;
wire      [7:0] n355;
wire      [7:0] n356;
wire      [7:0] n357;
wire      [7:0] n358;
wire      [7:0] n359;
wire      [7:0] n360;
wire      [7:0] n361;
wire      [7:0] n362;
wire      [7:0] n363;
wire      [7:0] n364;
wire      [7:0] n365;
wire      [7:0] n366;
wire      [7:0] n367;
wire      [7:0] n368;
wire      [7:0] n369;
wire      [7:0] n370;
wire      [7:0] n371;
wire      [7:0] n372;
wire      [7:0] n373;
wire      [7:0] n374;
wire      [7:0] n375;
wire      [7:0] n376;
wire      [7:0] n377;
wire      [7:0] n378;
wire      [7:0] n379;
wire      [7:0] n380;
wire      [7:0] n381;
wire      [7:0] n382;
wire      [7:0] n383;
wire      [7:0] n384;
wire      [7:0] n385;
wire      [7:0] n386;
wire      [7:0] n387;
wire      [7:0] n388;
wire      [7:0] n389;
wire      [7:0] n390;
wire      [7:0] n391;
wire      [7:0] n392;
wire      [7:0] n393;
wire      [7:0] n394;
wire      [7:0] n395;
wire     [15:0] n396;
wire     [23:0] n397;
wire     [31:0] n398;
wire     [39:0] n399;
wire     [47:0] n400;
wire     [55:0] n401;
wire     [63:0] n402;
wire     [71:0] n403;
wire     [71:0] n404;
wire     [71:0] n405;
wire     [71:0] n406;
wire     [71:0] n407;
wire     [71:0] n408;
wire     [71:0] n409;
wire     [71:0] n410;
wire     [71:0] n411;
wire     [71:0] n412;
wire     [71:0] n413;
wire     [71:0] n414;
wire     [71:0] n415;
wire     [71:0] n416;
wire     [71:0] n417;
wire            n418;
wire            n419;
wire            n420;
wire            n421;
wire            n422;
wire            n423;
wire            n424;
wire            n425;
wire            n426;
wire            n427;
wire            n428;
wire            n429;
wire            n430;
wire            n431;
wire            n432;
wire            n433;
wire            n434;
wire            n435;
wire      [7:0] n436;
wire      [7:0] n437;
wire      [7:0] n438;
wire      [7:0] n439;
wire      [7:0] n440;
wire      [7:0] n441;
wire      [7:0] n442;
wire      [7:0] n443;
wire      [7:0] n444;
wire     [15:0] n445;
wire     [23:0] n446;
wire     [31:0] n447;
wire     [39:0] n448;
wire     [47:0] n449;
wire     [55:0] n450;
wire     [63:0] n451;
wire     [71:0] n452;
wire      [7:0] n453;
wire      [7:0] n454;
wire      [7:0] n455;
wire      [7:0] n456;
wire      [7:0] n457;
wire      [7:0] n458;
wire      [7:0] n459;
wire      [7:0] n460;
wire      [7:0] n461;
wire     [15:0] n462;
wire     [23:0] n463;
wire     [31:0] n464;
wire     [39:0] n465;
wire     [47:0] n466;
wire     [55:0] n467;
wire     [63:0] n468;
wire     [71:0] n469;
wire      [7:0] n470;
wire      [7:0] n471;
wire      [7:0] n472;
wire      [7:0] n473;
wire      [7:0] n474;
wire      [7:0] n475;
wire      [7:0] n476;
wire      [7:0] n477;
wire      [7:0] n478;
wire     [15:0] n479;
wire     [23:0] n480;
wire     [31:0] n481;
wire     [39:0] n482;
wire     [47:0] n483;
wire     [55:0] n484;
wire     [63:0] n485;
wire     [71:0] n486;
wire      [7:0] n487;
wire      [7:0] n488;
wire      [7:0] n489;
wire      [7:0] n490;
wire      [7:0] n491;
wire      [7:0] n492;
wire      [7:0] n493;
wire      [7:0] n494;
wire      [7:0] n495;
wire     [15:0] n496;
wire     [23:0] n497;
wire     [31:0] n498;
wire     [39:0] n499;
wire     [47:0] n500;
wire     [55:0] n501;
wire     [63:0] n502;
wire     [71:0] n503;
wire      [7:0] n504;
wire      [7:0] n505;
wire      [7:0] n506;
wire      [7:0] n507;
wire      [7:0] n508;
wire      [7:0] n509;
wire      [7:0] n510;
wire      [7:0] n511;
wire      [7:0] n512;
wire     [15:0] n513;
wire     [23:0] n514;
wire     [31:0] n515;
wire     [39:0] n516;
wire     [47:0] n517;
wire     [55:0] n518;
wire     [63:0] n519;
wire     [71:0] n520;
wire      [7:0] n521;
wire      [7:0] n522;
wire      [7:0] n523;
wire      [7:0] n524;
wire      [7:0] n525;
wire      [7:0] n526;
wire      [7:0] n527;
wire      [7:0] n528;
wire      [7:0] n529;
wire     [15:0] n530;
wire     [23:0] n531;
wire     [31:0] n532;
wire     [39:0] n533;
wire     [47:0] n534;
wire     [55:0] n535;
wire     [63:0] n536;
wire     [71:0] n537;
wire      [7:0] n538;
wire      [7:0] n539;
wire      [7:0] n540;
wire      [7:0] n541;
wire      [7:0] n542;
wire      [7:0] n543;
wire      [7:0] n544;
wire      [7:0] n545;
wire      [7:0] n546;
wire     [15:0] n547;
wire     [23:0] n548;
wire     [31:0] n549;
wire     [39:0] n550;
wire     [47:0] n551;
wire     [55:0] n552;
wire     [63:0] n553;
wire     [71:0] n554;
wire      [7:0] n555;
wire      [7:0] n556;
wire      [7:0] n557;
wire      [7:0] n558;
wire      [7:0] n559;
wire      [7:0] n560;
wire      [7:0] n561;
wire      [7:0] n562;
wire      [7:0] n563;
wire     [15:0] n564;
wire     [23:0] n565;
wire     [31:0] n566;
wire     [39:0] n567;
wire     [47:0] n568;
wire     [55:0] n569;
wire     [63:0] n570;
wire     [71:0] n571;
wire      [7:0] n572;
wire      [7:0] n573;
wire      [7:0] n574;
wire      [7:0] n575;
wire      [7:0] n576;
wire      [7:0] n577;
wire      [7:0] n578;
wire      [7:0] n579;
wire      [7:0] n580;
wire     [15:0] n581;
wire     [23:0] n582;
wire     [31:0] n583;
wire     [39:0] n584;
wire     [47:0] n585;
wire     [55:0] n586;
wire     [63:0] n587;
wire     [71:0] n588;
wire    [143:0] n589;
wire    [215:0] n590;
wire    [287:0] n591;
wire    [359:0] n592;
wire    [431:0] n593;
wire    [503:0] n594;
wire    [575:0] n595;
wire    [647:0] n596;
wire    [647:0] n597;
wire    [647:0] n598;
wire    [647:0] n599;
wire    [647:0] n600;
wire    [647:0] n601;
wire    [647:0] n602;
wire    [647:0] n603;
wire    [647:0] n604;
wire    [647:0] n605;
wire    [647:0] n606;
wire    [647:0] n607;
wire    [647:0] n608;
wire    [647:0] n609;
wire            n610;
wire            n611;
wire            n612;
wire            n613;
wire            n614;
wire            n615;
wire            n616;
wire            n617;
wire            n618;
wire            n619;
wire            n620;
wire            n621;
wire            n622;
wire            n623;
wire            n624;
wire            n625;
wire            n626;
wire            n627;
wire      [8:0] LB2D_proc_0_addr0;
wire      [7:0] LB2D_proc_0_data0;
wire            n628;
wire            n629;
wire            n630;
wire            n631;
wire            n632;
wire            n633;
wire            n634;
wire            n635;
wire            n636;
wire            n637;
wire            n638;
wire            n639;
wire            n640;
wire            n641;
wire            n642;
wire            n643;
wire            n644;
wire            n645;
wire            n646;
wire      [8:0] LB2D_proc_1_addr0;
wire      [7:0] LB2D_proc_1_data0;
wire            n647;
wire            n648;
wire            n649;
wire      [8:0] LB2D_proc_2_addr0;
wire      [7:0] LB2D_proc_2_data0;
wire            n650;
wire            n651;
wire            n652;
wire      [8:0] LB2D_proc_3_addr0;
wire      [7:0] LB2D_proc_3_data0;
wire            n653;
wire            n654;
wire            n655;
wire      [8:0] LB2D_proc_4_addr0;
wire      [7:0] LB2D_proc_4_data0;
wire            n656;
wire            n657;
wire            n658;
wire      [8:0] LB2D_proc_5_addr0;
wire      [7:0] LB2D_proc_5_data0;
wire            n659;
wire            n660;
wire            n661;
wire      [8:0] LB2D_proc_6_addr0;
wire      [7:0] LB2D_proc_6_data0;
wire            n662;
wire            n663;
wire            n664;
wire      [8:0] LB2D_proc_7_addr0;
wire      [7:0] LB2D_proc_7_data0;
wire            n665;
wire            n666;
wire            n667;
wire            n668;
reg      [7:0] LB2D_proc_0[511:0];
reg      [7:0] LB2D_proc_1[511:0];
reg      [7:0] LB2D_proc_2[511:0];
reg      [7:0] LB2D_proc_3[511:0];
reg      [7:0] LB2D_proc_4[511:0];
reg      [7:0] LB2D_proc_5[511:0];
reg      [7:0] LB2D_proc_6[511:0];
reg      [7:0] LB2D_proc_7[511:0];
wire clk;
wire rst;
wire step;
assign n0 =  ( arg_0_TREADY ) == ( 1'd1 )  ;
assign n1 =  ( arg_0_TVALID ) == ( 1'd1 )  ;
assign n2 =  ( n0 ) & ( n1 )  ;
assign n3 =  ( arg_1_TVALID ) == ( 1'd0 )  ;
assign n4 =  ( n2 ) & ( n3 )  ;
assign n5 =  ( arg_1_TREADY ) == ( 1'd1 )  ;
assign n6 =  ( arg_1_TVALID ) == ( 1'd1 )  ;
assign n7 =  ( n5 ) & ( n6 )  ;
assign n8 =  ( arg_0_TREADY ) == ( 1'd0 )  ;
assign n9 =  ( n7 ) & ( n8 )  ;
assign n10 =  ( arg_0_TVALID ) == ( 1'd0 )  ;
assign n11 =  ( gb_exit_it_1 ) == ( 1'd0 )  ;
assign n12 =  ( stencil_stream_empty ) == ( 1'd0 )  ;
assign n13 =  ( n11 ) & ( n12 )  ;
assign n14 =  ( gb_exit_it_1 ) == ( 1'd1 )  ;
assign n15 =  ( gb_exit_it_8 ) == ( 1'd0 )  ;
assign n16 =  ( n14 ) & ( n15 )  ;
assign n17 =  ( n13 ) | ( n16 )  ;
assign n18 =  ( n10 ) & ( n17 )  ;
assign n19 =  ( slice_stream_empty ) == ( 1'd0 )  ;
assign n20 =  ( LB2D_shift_x ) != ( 9'd488 )  ;
assign n21 =  ( n19 ) & ( n20 )  ;
assign n22 =  ( stencil_stream_full ) == ( 1'd0 )  ;
assign n23 =  ( LB2D_shift_x ) < ( 9'd8 )  ;
assign n24 =  ( n22 ) | ( n23 )  ;
assign n25 =  ( n21 ) & ( n24 )  ;
assign n26 =  ( arg_1_TREADY ) == ( 1'd0 )  ;
assign n27 =  ( in_stream_full ) == ( 1'd0 )  ;
assign n28 =  ( n26 ) & ( n27 )  ;
assign n29 =  ( LB1D_it_1 ) == ( 1'd1 )  ;
assign n30 =  ( n28 ) & ( n29 )  ;
assign n31 =  ( n30 ) ? ( arg_1_TDATA ) : ( LB1D_in ) ;
assign n32 =  ( n25 ) ? ( LB1D_in ) : ( n31 ) ;
assign n33 =  ( n25 ) ? ( LB1D_buff ) : ( n32 ) ;
assign n34 =  ( n18 ) ? ( LB1D_buff ) : ( n33 ) ;
assign n35 =  ( n9 ) ? ( LB1D_buff ) : ( n34 ) ;
assign n36 =  ( n4 ) ? ( LB1D_buff ) : ( n35 ) ;
assign n37 =  ( n18 ) ? ( LB1D_in ) : ( n31 ) ;
assign n38 =  ( n9 ) ? ( LB1D_in ) : ( n37 ) ;
assign n39 =  ( n4 ) ? ( LB1D_in ) : ( n38 ) ;
assign n40 =  ( LB1D_it_1 ) == ( 1'd0 )  ;
assign n41 =  ( n28 ) & ( n40 )  ;
assign n42 =  ( n41 ) ? ( 1'd1 ) : ( LB1D_it_1 ) ;
assign n43 =  ( in_stream_empty ) == ( 1'd0 )  ;
assign n44 =  ( LB2D_proc_x ) != ( 9'd488 )  ;
assign n45 =  ( n43 ) & ( n44 )  ;
assign n46 =  ( slice_stream_full ) == ( 1'd0 )  ;
assign n47 =  ( LB2D_proc_y ) < ( 10'd8 )  ;
assign n48 =  ( n46 ) | ( n47 )  ;
assign n49 =  ( n45 ) & ( n48 )  ;
assign n50 =  ( LB1D_p_cnt ) + ( 19'd1 )  ;
assign n51 =  ( 19'd316224 ) - ( 19'd1 )  ;
assign n52 =  ( LB1D_p_cnt ) == ( n51 )  ;
assign n53 =  ( n52 ) ? ( 19'd0 ) : ( n50 ) ;
assign n54 =  ( n30 ) ? ( n53 ) : ( LB1D_p_cnt ) ;
assign n55 =  ( n41 ) ? ( n50 ) : ( n54 ) ;
assign n56 =  ( n49 ) ? ( LB1D_p_cnt ) : ( n55 ) ;
assign n57 =  ( n25 ) ? ( LB1D_p_cnt ) : ( n56 ) ;
assign n58 =  ( n18 ) ? ( LB1D_p_cnt ) : ( n57 ) ;
assign n59 =  ( n9 ) ? ( LB1D_p_cnt ) : ( n58 ) ;
assign n60 =  ( n4 ) ? ( LB1D_p_cnt ) : ( n59 ) ;
assign n61 =  ( LB2D_proc_w ) < ( 64'd7 )  ;
assign n62 =  ( LB2D_proc_x ) < ( 9'd488 )  ;
assign n63 =  ( LB2D_proc_w ) + ( 64'd1 )  ;
assign n64 =  ( n62 ) ? ( LB2D_proc_w ) : ( n63 ) ;
assign n65 =  ( n61 ) ? ( n64 ) : ( 64'd0 ) ;
assign n66 =  ( n30 ) ? ( LB2D_proc_w ) : ( LB2D_proc_w ) ;
assign n67 =  ( n49 ) ? ( n65 ) : ( n66 ) ;
assign n68 =  ( n25 ) ? ( LB2D_proc_w ) : ( n67 ) ;
assign n69 =  ( n18 ) ? ( LB2D_proc_w ) : ( n68 ) ;
assign n70 =  ( n9 ) ? ( LB2D_proc_w ) : ( n69 ) ;
assign n71 =  ( n4 ) ? ( LB2D_proc_w ) : ( n70 ) ;
assign n72 =  ( LB2D_proc_x ) == ( 9'd488 )  ;
assign n73 =  ( n43 ) & ( n72 )  ;
assign n74 =  ( n73 ) & ( n48 )  ;
assign n75 =  ( LB2D_proc_x ) + ( 9'd1 )  ;
assign n76 =  ( n30 ) ? ( LB2D_proc_x ) : ( LB2D_proc_x ) ;
assign n77 =  ( n49 ) ? ( n75 ) : ( n76 ) ;
assign n78 =  ( n74 ) ? ( 9'd0 ) : ( n77 ) ;
assign n79 =  ( n25 ) ? ( LB2D_proc_x ) : ( n78 ) ;
assign n80 =  ( n18 ) ? ( LB2D_proc_x ) : ( n79 ) ;
assign n81 =  ( n9 ) ? ( LB2D_proc_x ) : ( n80 ) ;
assign n82 =  ( n4 ) ? ( LB2D_proc_x ) : ( n81 ) ;
assign n83 =  ( LB2D_proc_y ) < ( 10'd488 )  ;
assign n84 =  ( n83 ) ? ( LB2D_proc_y ) : ( 10'd488 ) ;
assign n85 =  ( n30 ) ? ( LB2D_proc_y ) : ( LB2D_proc_y ) ;
assign n86 =  ( n49 ) ? ( n84 ) : ( n85 ) ;
assign n87 =  ( n25 ) ? ( LB2D_proc_y ) : ( n86 ) ;
assign n88 =  ( n18 ) ? ( LB2D_proc_y ) : ( n87 ) ;
assign n89 =  ( n9 ) ? ( LB2D_proc_y ) : ( n88 ) ;
assign n90 =  ( n4 ) ? ( LB2D_proc_y ) : ( n89 ) ;
assign n91 =  ( slice_stream_full ) == ( 1'd1 )  ;
assign n92 =  ( n91 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n93 =  ( n30 ) ? ( LB2D_shift_0 ) : ( LB2D_shift_0 ) ;
assign n94 =  ( n49 ) ? ( LB2D_shift_0 ) : ( n93 ) ;
assign n95 =  ( n25 ) ? ( n92 ) : ( n94 ) ;
assign n96 =  ( n18 ) ? ( LB2D_shift_0 ) : ( n95 ) ;
assign n97 =  ( n9 ) ? ( LB2D_shift_0 ) : ( n96 ) ;
assign n98 =  ( n4 ) ? ( LB2D_shift_0 ) : ( n97 ) ;
assign n99 =  ( n30 ) ? ( LB2D_shift_1 ) : ( LB2D_shift_1 ) ;
assign n100 =  ( n49 ) ? ( LB2D_shift_1 ) : ( n99 ) ;
assign n101 =  ( n25 ) ? ( LB2D_shift_0 ) : ( n100 ) ;
assign n102 =  ( n18 ) ? ( LB2D_shift_1 ) : ( n101 ) ;
assign n103 =  ( n9 ) ? ( LB2D_shift_1 ) : ( n102 ) ;
assign n104 =  ( n4 ) ? ( LB2D_shift_1 ) : ( n103 ) ;
assign n105 =  ( n30 ) ? ( LB2D_shift_2 ) : ( LB2D_shift_2 ) ;
assign n106 =  ( n49 ) ? ( LB2D_shift_2 ) : ( n105 ) ;
assign n107 =  ( n25 ) ? ( LB2D_shift_1 ) : ( n106 ) ;
assign n108 =  ( n18 ) ? ( LB2D_shift_2 ) : ( n107 ) ;
assign n109 =  ( n9 ) ? ( LB2D_shift_2 ) : ( n108 ) ;
assign n110 =  ( n4 ) ? ( LB2D_shift_2 ) : ( n109 ) ;
assign n111 =  ( n30 ) ? ( LB2D_shift_3 ) : ( LB2D_shift_3 ) ;
assign n112 =  ( n49 ) ? ( LB2D_shift_3 ) : ( n111 ) ;
assign n113 =  ( n25 ) ? ( LB2D_shift_2 ) : ( n112 ) ;
assign n114 =  ( n18 ) ? ( LB2D_shift_3 ) : ( n113 ) ;
assign n115 =  ( n9 ) ? ( LB2D_shift_3 ) : ( n114 ) ;
assign n116 =  ( n4 ) ? ( LB2D_shift_3 ) : ( n115 ) ;
assign n117 =  ( n30 ) ? ( LB2D_shift_4 ) : ( LB2D_shift_4 ) ;
assign n118 =  ( n49 ) ? ( LB2D_shift_4 ) : ( n117 ) ;
assign n119 =  ( n25 ) ? ( LB2D_shift_3 ) : ( n118 ) ;
assign n120 =  ( n18 ) ? ( LB2D_shift_4 ) : ( n119 ) ;
assign n121 =  ( n9 ) ? ( LB2D_shift_4 ) : ( n120 ) ;
assign n122 =  ( n4 ) ? ( LB2D_shift_4 ) : ( n121 ) ;
assign n123 =  ( n30 ) ? ( LB2D_shift_5 ) : ( LB2D_shift_5 ) ;
assign n124 =  ( n49 ) ? ( LB2D_shift_5 ) : ( n123 ) ;
assign n125 =  ( n25 ) ? ( LB2D_shift_4 ) : ( n124 ) ;
assign n126 =  ( n18 ) ? ( LB2D_shift_5 ) : ( n125 ) ;
assign n127 =  ( n9 ) ? ( LB2D_shift_5 ) : ( n126 ) ;
assign n128 =  ( n4 ) ? ( LB2D_shift_5 ) : ( n127 ) ;
assign n129 =  ( n30 ) ? ( LB2D_shift_6 ) : ( LB2D_shift_6 ) ;
assign n130 =  ( n49 ) ? ( LB2D_shift_6 ) : ( n129 ) ;
assign n131 =  ( n25 ) ? ( LB2D_shift_5 ) : ( n130 ) ;
assign n132 =  ( n18 ) ? ( LB2D_shift_6 ) : ( n131 ) ;
assign n133 =  ( n9 ) ? ( LB2D_shift_6 ) : ( n132 ) ;
assign n134 =  ( n4 ) ? ( LB2D_shift_6 ) : ( n133 ) ;
assign n135 =  ( n30 ) ? ( LB2D_shift_7 ) : ( LB2D_shift_7 ) ;
assign n136 =  ( n49 ) ? ( LB2D_shift_7 ) : ( n135 ) ;
assign n137 =  ( n25 ) ? ( LB2D_shift_6 ) : ( n136 ) ;
assign n138 =  ( n18 ) ? ( LB2D_shift_7 ) : ( n137 ) ;
assign n139 =  ( n9 ) ? ( LB2D_shift_7 ) : ( n138 ) ;
assign n140 =  ( n4 ) ? ( LB2D_shift_7 ) : ( n139 ) ;
assign n141 =  ( LB2D_shift_x ) + ( 9'd1 )  ;
assign n142 =  ( n30 ) ? ( LB2D_shift_x ) : ( LB2D_shift_x ) ;
assign n143 =  ( n49 ) ? ( LB2D_shift_x ) : ( n142 ) ;
assign n144 =  ( n25 ) ? ( n141 ) : ( n143 ) ;
assign n145 =  ( n18 ) ? ( LB2D_shift_x ) : ( n144 ) ;
assign n146 =  ( n9 ) ? ( LB2D_shift_x ) : ( n145 ) ;
assign n147 =  ( n4 ) ? ( LB2D_shift_x ) : ( n146 ) ;
assign n148 =  ( LB2D_shift_y ) < ( 10'd480 )  ;
assign n149 =  ( LB2D_shift_x ) < ( 9'd488 )  ;
assign n150 =  ( LB2D_shift_y ) + ( 10'd1 )  ;
assign n151 =  ( n149 ) ? ( LB2D_shift_y ) : ( n150 ) ;
assign n152 =  ( n148 ) ? ( n151 ) : ( 10'd480 ) ;
assign n153 =  ( n30 ) ? ( LB2D_shift_y ) : ( LB2D_shift_y ) ;
assign n154 =  ( n49 ) ? ( LB2D_shift_y ) : ( n153 ) ;
assign n155 =  ( n25 ) ? ( n152 ) : ( n154 ) ;
assign n156 =  ( n18 ) ? ( LB2D_shift_y ) : ( n155 ) ;
assign n157 =  ( n9 ) ? ( LB2D_shift_y ) : ( n156 ) ;
assign n158 =  ( n4 ) ? ( LB2D_shift_y ) : ( n157 ) ;
assign n159 =  ( stencil_stream_full ) == ( 1'd1 )  ;
assign n160 =  ( n159 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_0 ) ;
//assign n161 = gb_fun(n160) ;
gb_fun gb_fun_U (
        .stencil (n160),
        .result (n161)
        );

assign n162 =  ( n30 ) ? ( arg_0_TDATA ) : ( arg_0_TDATA ) ;
assign n163 =  ( n49 ) ? ( arg_0_TDATA ) : ( n162 ) ;
assign n164 =  ( n25 ) ? ( arg_0_TDATA ) : ( n163 ) ;
assign n165 =  ( n18 ) ? ( n161 ) : ( n164 ) ;
assign n166 =  ( n9 ) ? ( arg_0_TDATA ) : ( n165 ) ;
assign n167 =  ( n4 ) ? ( arg_0_TDATA ) : ( n166 ) ;
assign n168 =  ( gb_pp_it_8 ) == ( 1'd1 )  ;
assign n169 =  ( n168 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n170 =  ( n30 ) ? ( arg_0_TVALID ) : ( arg_0_TVALID ) ;
assign n171 =  ( n49 ) ? ( arg_0_TVALID ) : ( n170 ) ;
assign n172 =  ( n25 ) ? ( arg_0_TVALID ) : ( n171 ) ;
assign n173 =  ( n18 ) ? ( n169 ) : ( n172 ) ;
assign n174 =  ( n9 ) ? ( arg_0_TVALID ) : ( n173 ) ;
assign n175 =  ( n4 ) ? ( 1'd0 ) : ( n174 ) ;
assign n176 =  ( n30 ) ? ( 1'd1 ) : ( arg_1_TREADY ) ;
assign n177 =  ( n41 ) ? ( 1'd1 ) : ( n176 ) ;
assign n178 =  ( n49 ) ? ( arg_1_TREADY ) : ( n177 ) ;
assign n179 =  ( n25 ) ? ( arg_1_TREADY ) : ( n178 ) ;
assign n180 =  ( n18 ) ? ( arg_1_TREADY ) : ( n179 ) ;
assign n181 =  ( n9 ) ? ( 1'd0 ) : ( n180 ) ;
assign n182 =  ( n4 ) ? ( 1'd0 ) : ( n181 ) ;
assign n183 =  ( gb_p_cnt ) + ( 19'd1 )  ;
assign n184 =  ( n183 ) == ( 19'd307200 )  ;
assign n185 =  ( n184 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n186 =  ( n30 ) ? ( gb_exit_it_1 ) : ( gb_exit_it_1 ) ;
assign n187 =  ( n49 ) ? ( gb_exit_it_1 ) : ( n186 ) ;
assign n188 =  ( n25 ) ? ( gb_exit_it_1 ) : ( n187 ) ;
assign n189 =  ( n18 ) ? ( n185 ) : ( n188 ) ;
assign n190 =  ( n9 ) ? ( gb_exit_it_1 ) : ( n189 ) ;
assign n191 =  ( n4 ) ? ( gb_exit_it_1 ) : ( n190 ) ;
assign n192 =  ( n30 ) ? ( gb_exit_it_2 ) : ( gb_exit_it_2 ) ;
assign n193 =  ( n49 ) ? ( gb_exit_it_2 ) : ( n192 ) ;
assign n194 =  ( n25 ) ? ( gb_exit_it_2 ) : ( n193 ) ;
assign n195 =  ( n18 ) ? ( gb_exit_it_1 ) : ( n194 ) ;
assign n196 =  ( n9 ) ? ( gb_exit_it_2 ) : ( n195 ) ;
assign n197 =  ( n4 ) ? ( gb_exit_it_2 ) : ( n196 ) ;
assign n198 =  ( n30 ) ? ( gb_exit_it_3 ) : ( gb_exit_it_3 ) ;
assign n199 =  ( n49 ) ? ( gb_exit_it_3 ) : ( n198 ) ;
assign n200 =  ( n25 ) ? ( gb_exit_it_3 ) : ( n199 ) ;
assign n201 =  ( n18 ) ? ( gb_exit_it_2 ) : ( n200 ) ;
assign n202 =  ( n9 ) ? ( gb_exit_it_3 ) : ( n201 ) ;
assign n203 =  ( n4 ) ? ( gb_exit_it_3 ) : ( n202 ) ;
assign n204 =  ( n30 ) ? ( gb_exit_it_4 ) : ( gb_exit_it_4 ) ;
assign n205 =  ( n49 ) ? ( gb_exit_it_4 ) : ( n204 ) ;
assign n206 =  ( n25 ) ? ( gb_exit_it_4 ) : ( n205 ) ;
assign n207 =  ( n18 ) ? ( gb_exit_it_3 ) : ( n206 ) ;
assign n208 =  ( n9 ) ? ( gb_exit_it_4 ) : ( n207 ) ;
assign n209 =  ( n4 ) ? ( gb_exit_it_4 ) : ( n208 ) ;
assign n210 =  ( n30 ) ? ( gb_exit_it_5 ) : ( gb_exit_it_5 ) ;
assign n211 =  ( n49 ) ? ( gb_exit_it_5 ) : ( n210 ) ;
assign n212 =  ( n25 ) ? ( gb_exit_it_5 ) : ( n211 ) ;
assign n213 =  ( n18 ) ? ( gb_exit_it_4 ) : ( n212 ) ;
assign n214 =  ( n9 ) ? ( gb_exit_it_5 ) : ( n213 ) ;
assign n215 =  ( n4 ) ? ( gb_exit_it_5 ) : ( n214 ) ;
assign n216 =  ( n30 ) ? ( gb_exit_it_6 ) : ( gb_exit_it_6 ) ;
assign n217 =  ( n49 ) ? ( gb_exit_it_6 ) : ( n216 ) ;
assign n218 =  ( n25 ) ? ( gb_exit_it_6 ) : ( n217 ) ;
assign n219 =  ( n18 ) ? ( gb_exit_it_5 ) : ( n218 ) ;
assign n220 =  ( n9 ) ? ( gb_exit_it_6 ) : ( n219 ) ;
assign n221 =  ( n4 ) ? ( gb_exit_it_6 ) : ( n220 ) ;
assign n222 =  ( n30 ) ? ( gb_exit_it_7 ) : ( gb_exit_it_7 ) ;
assign n223 =  ( n49 ) ? ( gb_exit_it_7 ) : ( n222 ) ;
assign n224 =  ( n25 ) ? ( gb_exit_it_7 ) : ( n223 ) ;
assign n225 =  ( n18 ) ? ( gb_exit_it_6 ) : ( n224 ) ;
assign n226 =  ( n9 ) ? ( gb_exit_it_7 ) : ( n225 ) ;
assign n227 =  ( n4 ) ? ( gb_exit_it_7 ) : ( n226 ) ;
assign n228 =  ( n30 ) ? ( gb_exit_it_8 ) : ( gb_exit_it_8 ) ;
assign n229 =  ( n49 ) ? ( gb_exit_it_8 ) : ( n228 ) ;
assign n230 =  ( n25 ) ? ( gb_exit_it_8 ) : ( n229 ) ;
assign n231 =  ( n18 ) ? ( gb_exit_it_7 ) : ( n230 ) ;
assign n232 =  ( n9 ) ? ( gb_exit_it_8 ) : ( n231 ) ;
assign n233 =  ( n4 ) ? ( gb_exit_it_8 ) : ( n232 ) ;
assign n234 =  ( gb_p_cnt ) < ( 19'd307200 )  ;
assign n235 =  ( n234 ) ? ( n183 ) : ( 19'd307200 ) ;
assign n236 =  ( n30 ) ? ( gb_p_cnt ) : ( gb_p_cnt ) ;
assign n237 =  ( n49 ) ? ( gb_p_cnt ) : ( n236 ) ;
assign n238 =  ( n25 ) ? ( gb_p_cnt ) : ( n237 ) ;
assign n239 =  ( n18 ) ? ( n235 ) : ( n238 ) ;
assign n240 =  ( n9 ) ? ( gb_p_cnt ) : ( n239 ) ;
assign n241 =  ( n4 ) ? ( gb_p_cnt ) : ( n240 ) ;
assign n242 =  ( n30 ) ? ( gb_pp_it_1 ) : ( gb_pp_it_1 ) ;
assign n243 =  ( n49 ) ? ( gb_pp_it_1 ) : ( n242 ) ;
assign n244 =  ( n25 ) ? ( gb_pp_it_1 ) : ( n243 ) ;
assign n245 =  ( n18 ) ? ( 1'd1 ) : ( n244 ) ;
assign n246 =  ( n9 ) ? ( gb_pp_it_1 ) : ( n245 ) ;
assign n247 =  ( n4 ) ? ( gb_pp_it_1 ) : ( n246 ) ;
assign n248 =  ( n30 ) ? ( gb_pp_it_2 ) : ( gb_pp_it_2 ) ;
assign n249 =  ( n49 ) ? ( gb_pp_it_2 ) : ( n248 ) ;
assign n250 =  ( n25 ) ? ( gb_pp_it_2 ) : ( n249 ) ;
assign n251 =  ( n18 ) ? ( gb_pp_it_1 ) : ( n250 ) ;
assign n252 =  ( n9 ) ? ( gb_pp_it_2 ) : ( n251 ) ;
assign n253 =  ( n4 ) ? ( gb_pp_it_2 ) : ( n252 ) ;
assign n254 =  ( n30 ) ? ( gb_pp_it_3 ) : ( gb_pp_it_3 ) ;
assign n255 =  ( n49 ) ? ( gb_pp_it_3 ) : ( n254 ) ;
assign n256 =  ( n25 ) ? ( gb_pp_it_3 ) : ( n255 ) ;
assign n257 =  ( n18 ) ? ( gb_pp_it_2 ) : ( n256 ) ;
assign n258 =  ( n9 ) ? ( gb_pp_it_3 ) : ( n257 ) ;
assign n259 =  ( n4 ) ? ( gb_pp_it_3 ) : ( n258 ) ;
assign n260 =  ( n30 ) ? ( gb_pp_it_4 ) : ( gb_pp_it_4 ) ;
assign n261 =  ( n49 ) ? ( gb_pp_it_4 ) : ( n260 ) ;
assign n262 =  ( n25 ) ? ( gb_pp_it_4 ) : ( n261 ) ;
assign n263 =  ( n18 ) ? ( gb_pp_it_3 ) : ( n262 ) ;
assign n264 =  ( n9 ) ? ( gb_pp_it_4 ) : ( n263 ) ;
assign n265 =  ( n4 ) ? ( gb_pp_it_4 ) : ( n264 ) ;
assign n266 =  ( n30 ) ? ( gb_pp_it_5 ) : ( gb_pp_it_5 ) ;
assign n267 =  ( n49 ) ? ( gb_pp_it_5 ) : ( n266 ) ;
assign n268 =  ( n25 ) ? ( gb_pp_it_5 ) : ( n267 ) ;
assign n269 =  ( n18 ) ? ( gb_pp_it_4 ) : ( n268 ) ;
assign n270 =  ( n9 ) ? ( gb_pp_it_5 ) : ( n269 ) ;
assign n271 =  ( n4 ) ? ( gb_pp_it_5 ) : ( n270 ) ;
assign n272 =  ( n30 ) ? ( gb_pp_it_6 ) : ( gb_pp_it_6 ) ;
assign n273 =  ( n49 ) ? ( gb_pp_it_6 ) : ( n272 ) ;
assign n274 =  ( n25 ) ? ( gb_pp_it_6 ) : ( n273 ) ;
assign n275 =  ( n18 ) ? ( gb_pp_it_5 ) : ( n274 ) ;
assign n276 =  ( n9 ) ? ( gb_pp_it_6 ) : ( n275 ) ;
assign n277 =  ( n4 ) ? ( gb_pp_it_6 ) : ( n276 ) ;
assign n278 =  ( n30 ) ? ( gb_pp_it_7 ) : ( gb_pp_it_7 ) ;
assign n279 =  ( n49 ) ? ( gb_pp_it_7 ) : ( n278 ) ;
assign n280 =  ( n25 ) ? ( gb_pp_it_7 ) : ( n279 ) ;
assign n281 =  ( n18 ) ? ( gb_pp_it_6 ) : ( n280 ) ;
assign n282 =  ( n9 ) ? ( gb_pp_it_7 ) : ( n281 ) ;
assign n283 =  ( n4 ) ? ( gb_pp_it_7 ) : ( n282 ) ;
assign n284 =  ( n30 ) ? ( gb_pp_it_8 ) : ( gb_pp_it_8 ) ;
assign n285 =  ( n49 ) ? ( gb_pp_it_8 ) : ( n284 ) ;
assign n286 =  ( n25 ) ? ( gb_pp_it_8 ) : ( n285 ) ;
assign n287 =  ( n18 ) ? ( gb_pp_it_7 ) : ( n286 ) ;
assign n288 =  ( n9 ) ? ( gb_pp_it_8 ) : ( n287 ) ;
assign n289 =  ( n4 ) ? ( gb_pp_it_8 ) : ( n288 ) ;
assign n290 =  ( n30 ) ? ( gb_pp_it_9 ) : ( gb_pp_it_9 ) ;
assign n291 =  ( n49 ) ? ( gb_pp_it_9 ) : ( n290 ) ;
assign n292 =  ( n25 ) ? ( gb_pp_it_9 ) : ( n291 ) ;
assign n293 =  ( n18 ) ? ( gb_pp_it_8 ) : ( n292 ) ;
assign n294 =  ( n9 ) ? ( gb_pp_it_9 ) : ( n293 ) ;
assign n295 =  ( n4 ) ? ( gb_pp_it_9 ) : ( n294 ) ;
assign n296 =  ( n30 ) ? ( LB1D_buff ) : ( in_stream_buff_0 ) ;
assign n297 =  ( n49 ) ? ( in_stream_buff_0 ) : ( n296 ) ;
assign n298 =  ( n25 ) ? ( in_stream_buff_0 ) : ( n297 ) ;
assign n299 =  ( n18 ) ? ( in_stream_buff_0 ) : ( n298 ) ;
assign n300 =  ( n9 ) ? ( in_stream_buff_0 ) : ( n299 ) ;
assign n301 =  ( n4 ) ? ( in_stream_buff_0 ) : ( n300 ) ;
assign n302 =  ( n30 ) ? ( in_stream_buff_0 ) : ( in_stream_buff_1 ) ;
assign n303 =  ( n49 ) ? ( in_stream_buff_1 ) : ( n302 ) ;
assign n304 =  ( n25 ) ? ( in_stream_buff_1 ) : ( n303 ) ;
assign n305 =  ( n18 ) ? ( in_stream_buff_1 ) : ( n304 ) ;
assign n306 =  ( n9 ) ? ( in_stream_buff_1 ) : ( n305 ) ;
assign n307 =  ( n4 ) ? ( in_stream_buff_1 ) : ( n306 ) ;
assign n308 =  ( in_stream_full ) == ( 1'd1 )  ;
assign n309 =  ( n308 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n310 =  ( n30 ) ? ( 1'd0 ) : ( in_stream_empty ) ;
assign n311 =  ( n49 ) ? ( n309 ) : ( n310 ) ;
assign n312 =  ( n25 ) ? ( in_stream_empty ) : ( n311 ) ;
assign n313 =  ( n18 ) ? ( in_stream_empty ) : ( n312 ) ;
assign n314 =  ( n9 ) ? ( in_stream_empty ) : ( n313 ) ;
assign n315 =  ( n4 ) ? ( in_stream_empty ) : ( n314 ) ;
assign n316 =  ( in_stream_empty ) == ( 1'd1 )  ;
assign n317 =  ( n316 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n318 =  ( n30 ) ? ( n317 ) : ( in_stream_full ) ;
assign n319 =  ( n49 ) ? ( 1'd0 ) : ( n318 ) ;
assign n320 =  ( n25 ) ? ( in_stream_full ) : ( n319 ) ;
assign n321 =  ( n18 ) ? ( in_stream_full ) : ( n320 ) ;
assign n322 =  ( n9 ) ? ( in_stream_full ) : ( n321 ) ;
assign n323 =  ( n4 ) ? ( in_stream_full ) : ( n322 ) ;
assign n324 =  ( n308 ) ? ( in_stream_buff_1 ) : ( in_stream_buff_0 ) ;
assign n325 =  ( LB2D_proc_w ) == ( 64'd0 )  ;
assign n326 =  (  LB2D_proc_7 [ LB2D_proc_x ] )  ;
assign n327 =  ( LB2D_proc_w ) == ( 64'd1 )  ;
assign n328 =  (  LB2D_proc_0 [ LB2D_proc_x ] )  ;
assign n329 =  ( LB2D_proc_w ) == ( 64'd2 )  ;
assign n330 =  (  LB2D_proc_1 [ LB2D_proc_x ] )  ;
assign n331 =  ( LB2D_proc_w ) == ( 64'd3 )  ;
assign n332 =  (  LB2D_proc_2 [ LB2D_proc_x ] )  ;
assign n333 =  ( LB2D_proc_w ) == ( 64'd4 )  ;
assign n334 =  (  LB2D_proc_3 [ LB2D_proc_x ] )  ;
assign n335 =  ( LB2D_proc_w ) == ( 64'd5 )  ;
assign n336 =  (  LB2D_proc_4 [ LB2D_proc_x ] )  ;
assign n337 =  ( LB2D_proc_w ) == ( 64'd6 )  ;
assign n338 =  (  LB2D_proc_5 [ LB2D_proc_x ] )  ;
assign n339 =  (  LB2D_proc_6 [ LB2D_proc_x ] )  ;
assign n340 =  ( n337 ) ? ( n338 ) : ( n339 ) ;
assign n341 =  ( n335 ) ? ( n336 ) : ( n340 ) ;
assign n342 =  ( n333 ) ? ( n334 ) : ( n341 ) ;
assign n343 =  ( n331 ) ? ( n332 ) : ( n342 ) ;
assign n344 =  ( n329 ) ? ( n330 ) : ( n343 ) ;
assign n345 =  ( n327 ) ? ( n328 ) : ( n344 ) ;
assign n346 =  ( n325 ) ? ( n326 ) : ( n345 ) ;
assign n347 =  ( n337 ) ? ( n336 ) : ( n338 ) ;
assign n348 =  ( n335 ) ? ( n334 ) : ( n347 ) ;
assign n349 =  ( n333 ) ? ( n332 ) : ( n348 ) ;
assign n350 =  ( n331 ) ? ( n330 ) : ( n349 ) ;
assign n351 =  ( n329 ) ? ( n328 ) : ( n350 ) ;
assign n352 =  ( n327 ) ? ( n326 ) : ( n351 ) ;
assign n353 =  ( n325 ) ? ( n339 ) : ( n352 ) ;
assign n354 =  ( n337 ) ? ( n334 ) : ( n336 ) ;
assign n355 =  ( n335 ) ? ( n332 ) : ( n354 ) ;
assign n356 =  ( n333 ) ? ( n330 ) : ( n355 ) ;
assign n357 =  ( n331 ) ? ( n328 ) : ( n356 ) ;
assign n358 =  ( n329 ) ? ( n326 ) : ( n357 ) ;
assign n359 =  ( n327 ) ? ( n339 ) : ( n358 ) ;
assign n360 =  ( n325 ) ? ( n338 ) : ( n359 ) ;
assign n361 =  ( n337 ) ? ( n332 ) : ( n334 ) ;
assign n362 =  ( n335 ) ? ( n330 ) : ( n361 ) ;
assign n363 =  ( n333 ) ? ( n328 ) : ( n362 ) ;
assign n364 =  ( n331 ) ? ( n326 ) : ( n363 ) ;
assign n365 =  ( n329 ) ? ( n339 ) : ( n364 ) ;
assign n366 =  ( n327 ) ? ( n338 ) : ( n365 ) ;
assign n367 =  ( n325 ) ? ( n336 ) : ( n366 ) ;
assign n368 =  ( n337 ) ? ( n330 ) : ( n332 ) ;
assign n369 =  ( n335 ) ? ( n328 ) : ( n368 ) ;
assign n370 =  ( n333 ) ? ( n326 ) : ( n369 ) ;
assign n371 =  ( n331 ) ? ( n339 ) : ( n370 ) ;
assign n372 =  ( n329 ) ? ( n338 ) : ( n371 ) ;
assign n373 =  ( n327 ) ? ( n336 ) : ( n372 ) ;
assign n374 =  ( n325 ) ? ( n334 ) : ( n373 ) ;
assign n375 =  ( n337 ) ? ( n328 ) : ( n330 ) ;
assign n376 =  ( n335 ) ? ( n326 ) : ( n375 ) ;
assign n377 =  ( n333 ) ? ( n339 ) : ( n376 ) ;
assign n378 =  ( n331 ) ? ( n338 ) : ( n377 ) ;
assign n379 =  ( n329 ) ? ( n336 ) : ( n378 ) ;
assign n380 =  ( n327 ) ? ( n334 ) : ( n379 ) ;
assign n381 =  ( n325 ) ? ( n332 ) : ( n380 ) ;
assign n382 =  ( n337 ) ? ( n326 ) : ( n328 ) ;
assign n383 =  ( n335 ) ? ( n339 ) : ( n382 ) ;
assign n384 =  ( n333 ) ? ( n338 ) : ( n383 ) ;
assign n385 =  ( n331 ) ? ( n336 ) : ( n384 ) ;
assign n386 =  ( n329 ) ? ( n334 ) : ( n385 ) ;
assign n387 =  ( n327 ) ? ( n332 ) : ( n386 ) ;
assign n388 =  ( n325 ) ? ( n330 ) : ( n387 ) ;
assign n389 =  ( n337 ) ? ( n339 ) : ( n326 ) ;
assign n390 =  ( n335 ) ? ( n338 ) : ( n389 ) ;
assign n391 =  ( n333 ) ? ( n336 ) : ( n390 ) ;
assign n392 =  ( n331 ) ? ( n334 ) : ( n391 ) ;
assign n393 =  ( n329 ) ? ( n332 ) : ( n392 ) ;
assign n394 =  ( n327 ) ? ( n330 ) : ( n393 ) ;
assign n395 =  ( n325 ) ? ( n328 ) : ( n394 ) ;
assign n396 =  { ( n388 ) , ( n395 ) }  ;
assign n397 =  { ( n381 ) , ( n396 ) }  ;
assign n398 =  { ( n374 ) , ( n397 ) }  ;
assign n399 =  { ( n367 ) , ( n398 ) }  ;
assign n400 =  { ( n360 ) , ( n399 ) }  ;
assign n401 =  { ( n353 ) , ( n400 ) }  ;
assign n402 =  { ( n346 ) , ( n401 ) }  ;
assign n403 =  { ( n324 ) , ( n402 ) }  ;
assign n404 =  ( n47 ) ? ( slice_stream_buff_0 ) : ( n403 ) ;
assign n405 =  ( n30 ) ? ( slice_stream_buff_0 ) : ( slice_stream_buff_0 ) ;
assign n406 =  ( n49 ) ? ( n404 ) : ( n405 ) ;
assign n407 =  ( n25 ) ? ( slice_stream_buff_0 ) : ( n406 ) ;
assign n408 =  ( n18 ) ? ( slice_stream_buff_0 ) : ( n407 ) ;
assign n409 =  ( n9 ) ? ( slice_stream_buff_0 ) : ( n408 ) ;
assign n410 =  ( n4 ) ? ( slice_stream_buff_0 ) : ( n409 ) ;
assign n411 =  ( n47 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n412 =  ( n30 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_1 ) ;
assign n413 =  ( n49 ) ? ( n411 ) : ( n412 ) ;
assign n414 =  ( n25 ) ? ( slice_stream_buff_1 ) : ( n413 ) ;
assign n415 =  ( n18 ) ? ( slice_stream_buff_1 ) : ( n414 ) ;
assign n416 =  ( n9 ) ? ( slice_stream_buff_1 ) : ( n415 ) ;
assign n417 =  ( n4 ) ? ( slice_stream_buff_1 ) : ( n416 ) ;
assign n418 =  ( n91 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n419 =  ( n47 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n420 =  ( n30 ) ? ( slice_stream_empty ) : ( slice_stream_empty ) ;
assign n421 =  ( n49 ) ? ( n419 ) : ( n420 ) ;
assign n422 =  ( n25 ) ? ( n418 ) : ( n421 ) ;
assign n423 =  ( n18 ) ? ( slice_stream_empty ) : ( n422 ) ;
assign n424 =  ( n9 ) ? ( slice_stream_empty ) : ( n423 ) ;
assign n425 =  ( n4 ) ? ( slice_stream_empty ) : ( n424 ) ;
assign n426 =  ( slice_stream_empty ) == ( 1'd1 )  ;
assign n427 =  ( n426 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n428 =  ( n47 ) ? ( 1'd0 ) : ( n427 ) ;
assign n429 =  ( n30 ) ? ( slice_stream_full ) : ( slice_stream_full ) ;
assign n430 =  ( n49 ) ? ( n428 ) : ( n429 ) ;
assign n431 =  ( n25 ) ? ( 1'd0 ) : ( n430 ) ;
assign n432 =  ( n18 ) ? ( slice_stream_full ) : ( n431 ) ;
assign n433 =  ( n9 ) ? ( slice_stream_full ) : ( n432 ) ;
assign n434 =  ( n4 ) ? ( slice_stream_full ) : ( n433 ) ;
assign n435 =  ( LB2D_shift_x ) >= ( 9'd8 )  ;
assign n436 = n92[71:64] ;
assign n437 = LB2D_shift_0[71:64] ;
assign n438 = LB2D_shift_1[71:64] ;
assign n439 = LB2D_shift_2[71:64] ;
assign n440 = LB2D_shift_3[71:64] ;
assign n441 = LB2D_shift_4[71:64] ;
assign n442 = LB2D_shift_5[71:64] ;
assign n443 = LB2D_shift_6[71:64] ;
assign n444 = LB2D_shift_7[71:64] ;
assign n445 =  { ( n443 ) , ( n444 ) }  ;
assign n446 =  { ( n442 ) , ( n445 ) }  ;
assign n447 =  { ( n441 ) , ( n446 ) }  ;
assign n448 =  { ( n440 ) , ( n447 ) }  ;
assign n449 =  { ( n439 ) , ( n448 ) }  ;
assign n450 =  { ( n438 ) , ( n449 ) }  ;
assign n451 =  { ( n437 ) , ( n450 ) }  ;
assign n452 =  { ( n436 ) , ( n451 ) }  ;
assign n453 = n92[63:56] ;
assign n454 = LB2D_shift_0[63:56] ;
assign n455 = LB2D_shift_1[63:56] ;
assign n456 = LB2D_shift_2[63:56] ;
assign n457 = LB2D_shift_3[63:56] ;
assign n458 = LB2D_shift_4[63:56] ;
assign n459 = LB2D_shift_5[63:56] ;
assign n460 = LB2D_shift_6[63:56] ;
assign n461 = LB2D_shift_7[63:56] ;
assign n462 =  { ( n460 ) , ( n461 ) }  ;
assign n463 =  { ( n459 ) , ( n462 ) }  ;
assign n464 =  { ( n458 ) , ( n463 ) }  ;
assign n465 =  { ( n457 ) , ( n464 ) }  ;
assign n466 =  { ( n456 ) , ( n465 ) }  ;
assign n467 =  { ( n455 ) , ( n466 ) }  ;
assign n468 =  { ( n454 ) , ( n467 ) }  ;
assign n469 =  { ( n453 ) , ( n468 ) }  ;
assign n470 = n92[55:48] ;
assign n471 = LB2D_shift_0[55:48] ;
assign n472 = LB2D_shift_1[55:48] ;
assign n473 = LB2D_shift_2[55:48] ;
assign n474 = LB2D_shift_3[55:48] ;
assign n475 = LB2D_shift_4[55:48] ;
assign n476 = LB2D_shift_5[55:48] ;
assign n477 = LB2D_shift_6[55:48] ;
assign n478 = LB2D_shift_7[55:48] ;
assign n479 =  { ( n477 ) , ( n478 ) }  ;
assign n480 =  { ( n476 ) , ( n479 ) }  ;
assign n481 =  { ( n475 ) , ( n480 ) }  ;
assign n482 =  { ( n474 ) , ( n481 ) }  ;
assign n483 =  { ( n473 ) , ( n482 ) }  ;
assign n484 =  { ( n472 ) , ( n483 ) }  ;
assign n485 =  { ( n471 ) , ( n484 ) }  ;
assign n486 =  { ( n470 ) , ( n485 ) }  ;
assign n487 = n92[47:40] ;
assign n488 = LB2D_shift_0[47:40] ;
assign n489 = LB2D_shift_1[47:40] ;
assign n490 = LB2D_shift_2[47:40] ;
assign n491 = LB2D_shift_3[47:40] ;
assign n492 = LB2D_shift_4[47:40] ;
assign n493 = LB2D_shift_5[47:40] ;
assign n494 = LB2D_shift_6[47:40] ;
assign n495 = LB2D_shift_7[47:40] ;
assign n496 =  { ( n494 ) , ( n495 ) }  ;
assign n497 =  { ( n493 ) , ( n496 ) }  ;
assign n498 =  { ( n492 ) , ( n497 ) }  ;
assign n499 =  { ( n491 ) , ( n498 ) }  ;
assign n500 =  { ( n490 ) , ( n499 ) }  ;
assign n501 =  { ( n489 ) , ( n500 ) }  ;
assign n502 =  { ( n488 ) , ( n501 ) }  ;
assign n503 =  { ( n487 ) , ( n502 ) }  ;
assign n504 = n92[39:32] ;
assign n505 = LB2D_shift_0[39:32] ;
assign n506 = LB2D_shift_1[39:32] ;
assign n507 = LB2D_shift_2[39:32] ;
assign n508 = LB2D_shift_3[39:32] ;
assign n509 = LB2D_shift_4[39:32] ;
assign n510 = LB2D_shift_5[39:32] ;
assign n511 = LB2D_shift_6[39:32] ;
assign n512 = LB2D_shift_7[39:32] ;
assign n513 =  { ( n511 ) , ( n512 ) }  ;
assign n514 =  { ( n510 ) , ( n513 ) }  ;
assign n515 =  { ( n509 ) , ( n514 ) }  ;
assign n516 =  { ( n508 ) , ( n515 ) }  ;
assign n517 =  { ( n507 ) , ( n516 ) }  ;
assign n518 =  { ( n506 ) , ( n517 ) }  ;
assign n519 =  { ( n505 ) , ( n518 ) }  ;
assign n520 =  { ( n504 ) , ( n519 ) }  ;
assign n521 = n92[31:24] ;
assign n522 = LB2D_shift_0[31:24] ;
assign n523 = LB2D_shift_1[31:24] ;
assign n524 = LB2D_shift_2[31:24] ;
assign n525 = LB2D_shift_3[31:24] ;
assign n526 = LB2D_shift_4[31:24] ;
assign n527 = LB2D_shift_5[31:24] ;
assign n528 = LB2D_shift_6[31:24] ;
assign n529 = LB2D_shift_7[31:24] ;
assign n530 =  { ( n528 ) , ( n529 ) }  ;
assign n531 =  { ( n527 ) , ( n530 ) }  ;
assign n532 =  { ( n526 ) , ( n531 ) }  ;
assign n533 =  { ( n525 ) , ( n532 ) }  ;
assign n534 =  { ( n524 ) , ( n533 ) }  ;
assign n535 =  { ( n523 ) , ( n534 ) }  ;
assign n536 =  { ( n522 ) , ( n535 ) }  ;
assign n537 =  { ( n521 ) , ( n536 ) }  ;
assign n538 = n92[23:16] ;
assign n539 = LB2D_shift_0[23:16] ;
assign n540 = LB2D_shift_1[23:16] ;
assign n541 = LB2D_shift_2[23:16] ;
assign n542 = LB2D_shift_3[23:16] ;
assign n543 = LB2D_shift_4[23:16] ;
assign n544 = LB2D_shift_5[23:16] ;
assign n545 = LB2D_shift_6[23:16] ;
assign n546 = LB2D_shift_7[23:16] ;
assign n547 =  { ( n545 ) , ( n546 ) }  ;
assign n548 =  { ( n544 ) , ( n547 ) }  ;
assign n549 =  { ( n543 ) , ( n548 ) }  ;
assign n550 =  { ( n542 ) , ( n549 ) }  ;
assign n551 =  { ( n541 ) , ( n550 ) }  ;
assign n552 =  { ( n540 ) , ( n551 ) }  ;
assign n553 =  { ( n539 ) , ( n552 ) }  ;
assign n554 =  { ( n538 ) , ( n553 ) }  ;
assign n555 = n92[15:8] ;
assign n556 = LB2D_shift_0[15:8] ;
assign n557 = LB2D_shift_1[15:8] ;
assign n558 = LB2D_shift_2[15:8] ;
assign n559 = LB2D_shift_3[15:8] ;
assign n560 = LB2D_shift_4[15:8] ;
assign n561 = LB2D_shift_5[15:8] ;
assign n562 = LB2D_shift_6[15:8] ;
assign n563 = LB2D_shift_7[15:8] ;
assign n564 =  { ( n562 ) , ( n563 ) }  ;
assign n565 =  { ( n561 ) , ( n564 ) }  ;
assign n566 =  { ( n560 ) , ( n565 ) }  ;
assign n567 =  { ( n559 ) , ( n566 ) }  ;
assign n568 =  { ( n558 ) , ( n567 ) }  ;
assign n569 =  { ( n557 ) , ( n568 ) }  ;
assign n570 =  { ( n556 ) , ( n569 ) }  ;
assign n571 =  { ( n555 ) , ( n570 ) }  ;
assign n572 = n92[7:0] ;
assign n573 = LB2D_shift_0[7:0] ;
assign n574 = LB2D_shift_1[7:0] ;
assign n575 = LB2D_shift_2[7:0] ;
assign n576 = LB2D_shift_3[7:0] ;
assign n577 = LB2D_shift_4[7:0] ;
assign n578 = LB2D_shift_5[7:0] ;
assign n579 = LB2D_shift_6[7:0] ;
assign n580 = LB2D_shift_7[7:0] ;
assign n581 =  { ( n579 ) , ( n580 ) }  ;
assign n582 =  { ( n578 ) , ( n581 ) }  ;
assign n583 =  { ( n577 ) , ( n582 ) }  ;
assign n584 =  { ( n576 ) , ( n583 ) }  ;
assign n585 =  { ( n575 ) , ( n584 ) }  ;
assign n586 =  { ( n574 ) , ( n585 ) }  ;
assign n587 =  { ( n573 ) , ( n586 ) }  ;
assign n588 =  { ( n572 ) , ( n587 ) }  ;
assign n589 =  { ( n571 ) , ( n588 ) }  ;
assign n590 =  { ( n554 ) , ( n589 ) }  ;
assign n591 =  { ( n537 ) , ( n590 ) }  ;
assign n592 =  { ( n520 ) , ( n591 ) }  ;
assign n593 =  { ( n503 ) , ( n592 ) }  ;
assign n594 =  { ( n486 ) , ( n593 ) }  ;
assign n595 =  { ( n469 ) , ( n594 ) }  ;
assign n596 =  { ( n452 ) , ( n595 ) }  ;
assign n597 =  ( n435 ) ? ( n596 ) : ( stencil_stream_buff_0 ) ;
assign n598 =  ( n30 ) ? ( stencil_stream_buff_0 ) : ( stencil_stream_buff_0 ) ;
assign n599 =  ( n49 ) ? ( stencil_stream_buff_0 ) : ( n598 ) ;
assign n600 =  ( n25 ) ? ( n597 ) : ( n599 ) ;
assign n601 =  ( n18 ) ? ( stencil_stream_buff_0 ) : ( n600 ) ;
assign n602 =  ( n9 ) ? ( stencil_stream_buff_0 ) : ( n601 ) ;
assign n603 =  ( n4 ) ? ( stencil_stream_buff_0 ) : ( n602 ) ;
assign n604 =  ( n30 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_1 ) ;
assign n605 =  ( n49 ) ? ( stencil_stream_buff_1 ) : ( n604 ) ;
assign n606 =  ( n25 ) ? ( stencil_stream_buff_0 ) : ( n605 ) ;
assign n607 =  ( n18 ) ? ( stencil_stream_buff_1 ) : ( n606 ) ;
assign n608 =  ( n9 ) ? ( stencil_stream_buff_1 ) : ( n607 ) ;
assign n609 =  ( n4 ) ? ( stencil_stream_buff_1 ) : ( n608 ) ;
assign n610 =  ( n159 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n611 =  ( n23 ) ? ( stencil_stream_empty ) : ( 1'd0 ) ;
assign n612 =  ( n30 ) ? ( stencil_stream_empty ) : ( stencil_stream_empty ) ;
assign n613 =  ( n49 ) ? ( stencil_stream_empty ) : ( n612 ) ;
assign n614 =  ( n25 ) ? ( n611 ) : ( n613 ) ;
assign n615 =  ( n18 ) ? ( n610 ) : ( n614 ) ;
assign n616 =  ( n9 ) ? ( stencil_stream_empty ) : ( n615 ) ;
assign n617 =  ( n4 ) ? ( stencil_stream_empty ) : ( n616 ) ;
assign n618 =  ( n14 ) ? ( 1'd0 ) : ( 1'd0 ) ;
assign n619 =  ( stencil_stream_empty ) == ( 1'd1 )  ;
assign n620 =  ( n619 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n621 =  ( n23 ) ? ( stencil_stream_full ) : ( n620 ) ;
assign n622 =  ( n30 ) ? ( stencil_stream_full ) : ( stencil_stream_full ) ;
assign n623 =  ( n49 ) ? ( stencil_stream_full ) : ( n622 ) ;
assign n624 =  ( n25 ) ? ( n621 ) : ( n623 ) ;
assign n625 =  ( n18 ) ? ( n618 ) : ( n624 ) ;
assign n626 =  ( n9 ) ? ( stencil_stream_full ) : ( n625 ) ;
assign n627 =  ( n4 ) ? ( stencil_stream_full ) : ( n626 ) ;
assign n628 = ~ ( n4 ) ;
assign n629 = ~ ( n9 ) ;
assign n630 =  ( n628 ) & ( n629 )  ;
assign n631 = ~ ( n18 ) ;
assign n632 =  ( n630 ) & ( n631 )  ;
assign n633 = ~ ( n25 ) ;
assign n634 =  ( n632 ) & ( n633 )  ;
assign n635 = ~ ( n49 ) ;
assign n636 =  ( n634 ) & ( n635 )  ;
assign n637 = ~ ( n30 ) ;
assign n638 =  ( n636 ) & ( n637 )  ;
assign n639 =  ( n636 ) & ( n30 )  ;
assign n640 =  ( n634 ) & ( n49 )  ;
assign n641 = ~ ( n325 ) ;
assign n642 =  ( n640 ) & ( n641 )  ;
assign n643 =  ( n640 ) & ( n325 )  ;
assign n644 =  ( n632 ) & ( n25 )  ;
assign n645 =  ( n630 ) & ( n18 )  ;
assign n646 =  ( n628 ) & ( n9 )  ;
assign LB2D_proc_0_addr0 = n643 ? (LB2D_proc_x) : (0);
assign LB2D_proc_0_data0 = n643 ? (n324) : (LB2D_proc_0[0]);
assign n647 = ~ ( n327 ) ;
assign n648 =  ( n640 ) & ( n647 )  ;
assign n649 =  ( n640 ) & ( n327 )  ;
assign LB2D_proc_1_addr0 = n649 ? (LB2D_proc_x) : (0);
assign LB2D_proc_1_data0 = n649 ? (n324) : (LB2D_proc_1[0]);
assign n650 = ~ ( n329 ) ;
assign n651 =  ( n640 ) & ( n650 )  ;
assign n652 =  ( n640 ) & ( n329 )  ;
assign LB2D_proc_2_addr0 = n652 ? (LB2D_proc_x) : (0);
assign LB2D_proc_2_data0 = n652 ? (n324) : (LB2D_proc_2[0]);
assign n653 = ~ ( n331 ) ;
assign n654 =  ( n640 ) & ( n653 )  ;
assign n655 =  ( n640 ) & ( n331 )  ;
assign LB2D_proc_3_addr0 = n655 ? (LB2D_proc_x) : (0);
assign LB2D_proc_3_data0 = n655 ? (n324) : (LB2D_proc_3[0]);
assign n656 = ~ ( n333 ) ;
assign n657 =  ( n640 ) & ( n656 )  ;
assign n658 =  ( n640 ) & ( n333 )  ;
assign LB2D_proc_4_addr0 = n658 ? (LB2D_proc_x) : (0);
assign LB2D_proc_4_data0 = n658 ? (n324) : (LB2D_proc_4[0]);
assign n659 = ~ ( n335 ) ;
assign n660 =  ( n640 ) & ( n659 )  ;
assign n661 =  ( n640 ) & ( n335 )  ;
assign LB2D_proc_5_addr0 = n661 ? (LB2D_proc_x) : (0);
assign LB2D_proc_5_data0 = n661 ? (n324) : (LB2D_proc_5[0]);
assign n662 = ~ ( n337 ) ;
assign n663 =  ( n640 ) & ( n662 )  ;
assign n664 =  ( n640 ) & ( n337 )  ;
assign LB2D_proc_6_addr0 = n664 ? (LB2D_proc_x) : (0);
assign LB2D_proc_6_data0 = n664 ? (n324) : (LB2D_proc_6[0]);
assign n665 =  ( LB2D_proc_w ) == ( 64'd7 )  ;
assign n666 = ~ ( n665 ) ;
assign n667 =  ( n640 ) & ( n666 )  ;
assign n668 =  ( n640 ) & ( n665 )  ;
assign LB2D_proc_7_addr0 = n668 ? (LB2D_proc_x) : (0);
assign LB2D_proc_7_data0 = n668 ? (n324) : (LB2D_proc_7[0]);
/*
function [7:0] gb_fun ;
input [647:0] arg0;
    begin
//TODO: Add the specific function HERE.    end
endfunction
*/

always @(posedge clk) begin
   if(rst) begin
       LB1D_buff <= LB1D_buff;
       LB1D_in <= LB1D_in;
       LB1D_it_1 <= LB1D_it_1;
       LB1D_p_cnt <= LB1D_p_cnt;
       LB2D_proc_w <= LB2D_proc_w;
       LB2D_proc_x <= LB2D_proc_x;
       LB2D_proc_y <= LB2D_proc_y;
       LB2D_shift_0 <= LB2D_shift_0;
       LB2D_shift_1 <= LB2D_shift_1;
       LB2D_shift_2 <= LB2D_shift_2;
       LB2D_shift_3 <= LB2D_shift_3;
       LB2D_shift_4 <= LB2D_shift_4;
       LB2D_shift_5 <= LB2D_shift_5;
       LB2D_shift_6 <= LB2D_shift_6;
       LB2D_shift_7 <= LB2D_shift_7;
       LB2D_shift_x <= LB2D_shift_x;
       LB2D_shift_y <= LB2D_shift_y;
       arg_0_TDATA <= arg_0_TDATA;
       arg_0_TVALID <= arg_0_TVALID;
       arg_1_TREADY <= arg_1_TREADY;
       gb_exit_it_1 <= gb_exit_it_1;
       gb_exit_it_2 <= gb_exit_it_2;
       gb_exit_it_3 <= gb_exit_it_3;
       gb_exit_it_4 <= gb_exit_it_4;
       gb_exit_it_5 <= gb_exit_it_5;
       gb_exit_it_6 <= gb_exit_it_6;
       gb_exit_it_7 <= gb_exit_it_7;
       gb_exit_it_8 <= gb_exit_it_8;
       gb_p_cnt <= gb_p_cnt;
       gb_pp_it_1 <= gb_pp_it_1;
       gb_pp_it_2 <= gb_pp_it_2;
       gb_pp_it_3 <= gb_pp_it_3;
       gb_pp_it_4 <= gb_pp_it_4;
       gb_pp_it_5 <= gb_pp_it_5;
       gb_pp_it_6 <= gb_pp_it_6;
       gb_pp_it_7 <= gb_pp_it_7;
       gb_pp_it_8 <= gb_pp_it_8;
       gb_pp_it_9 <= gb_pp_it_9;
       in_stream_buff_0 <= in_stream_buff_0;
       in_stream_buff_1 <= in_stream_buff_1;
       in_stream_empty <= in_stream_empty;
       in_stream_full <= in_stream_full;
       slice_stream_buff_0 <= slice_stream_buff_0;
       slice_stream_buff_1 <= slice_stream_buff_1;
       slice_stream_empty <= slice_stream_empty;
       slice_stream_full <= slice_stream_full;
       stencil_stream_buff_0 <= stencil_stream_buff_0;
       stencil_stream_buff_1 <= stencil_stream_buff_1;
       stencil_stream_empty <= stencil_stream_empty;
       stencil_stream_full <= stencil_stream_full;
   end
   else if(step) begin
       LB1D_buff <= n36;
       LB1D_in <= n39;
       LB1D_it_1 <= n42;
       LB1D_p_cnt <= n60;
       LB2D_proc_w <= n71;
       LB2D_proc_x <= n82;
       LB2D_proc_y <= n90;
       LB2D_shift_0 <= n98;
       LB2D_shift_1 <= n104;
       LB2D_shift_2 <= n110;
       LB2D_shift_3 <= n116;
       LB2D_shift_4 <= n122;
       LB2D_shift_5 <= n128;
       LB2D_shift_6 <= n134;
       LB2D_shift_7 <= n140;
       LB2D_shift_x <= n147;
       LB2D_shift_y <= n158;
       arg_0_TDATA <= n167;
       arg_0_TVALID <= n175;
       arg_1_TREADY <= n182;
       gb_exit_it_1 <= n191;
       gb_exit_it_2 <= n197;
       gb_exit_it_3 <= n203;
       gb_exit_it_4 <= n209;
       gb_exit_it_5 <= n215;
       gb_exit_it_6 <= n221;
       gb_exit_it_7 <= n227;
       gb_exit_it_8 <= n233;
       gb_p_cnt <= n241;
       gb_pp_it_1 <= n247;
       gb_pp_it_2 <= n253;
       gb_pp_it_3 <= n259;
       gb_pp_it_4 <= n265;
       gb_pp_it_5 <= n271;
       gb_pp_it_6 <= n277;
       gb_pp_it_7 <= n283;
       gb_pp_it_8 <= n289;
       gb_pp_it_9 <= n295;
       in_stream_buff_0 <= n301;
       in_stream_buff_1 <= n307;
       in_stream_empty <= n315;
       in_stream_full <= n323;
       slice_stream_buff_0 <= n410;
       slice_stream_buff_1 <= n417;
       slice_stream_empty <= n425;
       slice_stream_full <= n434;
       stencil_stream_buff_0 <= n603;
       stencil_stream_buff_1 <= n609;
       stencil_stream_empty <= n617;
       stencil_stream_full <= n627;
       LB2D_proc_0 [ LB2D_proc_0_addr0 ] <= LB2D_proc_0_data0;
       LB2D_proc_1 [ LB2D_proc_1_addr0 ] <= LB2D_proc_1_data0;
       LB2D_proc_2 [ LB2D_proc_2_addr0 ] <= LB2D_proc_2_data0;
       LB2D_proc_3 [ LB2D_proc_3_addr0 ] <= LB2D_proc_3_data0;
       LB2D_proc_4 [ LB2D_proc_4_addr0 ] <= LB2D_proc_4_data0;
       LB2D_proc_5 [ LB2D_proc_5_addr0 ] <= LB2D_proc_5_data0;
       LB2D_proc_6 [ LB2D_proc_6_addr0 ] <= LB2D_proc_6_data0;
       LB2D_proc_7 [ LB2D_proc_7_addr0 ] <= LB2D_proc_7_data0;
   end
end
endmodule
