module GB(
arg_0_TREADY,
arg_1_TDATA,
arg_1_TVALID,
RAM_w,
RAM_x,
RAM_y,
arg_0_TDATA,
arg_0_TVALID,
arg_1_TREADY,
proc_in,
stencil_0,
stencil_1,
stencil_2,
stencil_3,
stencil_4,
stencil_5,
stencil_6,
stencil_7,
stencil_8,
clk,rst,
step
);
input            arg_0_TREADY;
input      [7:0] arg_1_TDATA;
input            arg_1_TVALID;
input clk;
input rst;
input step;
output      [2:0] RAM_w;
output      [8:0] RAM_x;
output      [9:0] RAM_y;
output      [7:0] arg_0_TDATA;
output            arg_0_TVALID;
output            arg_1_TREADY;
output    [647:0] proc_in;
output     [71:0] stencil_0;
output     [71:0] stencil_1;
output     [71:0] stencil_2;
output     [71:0] stencil_3;
output     [71:0] stencil_4;
output     [71:0] stencil_5;
output     [71:0] stencil_6;
output     [71:0] stencil_7;
output     [71:0] stencil_8;
reg      [2:0] RAM_w;
reg      [8:0] RAM_x;
reg      [9:0] RAM_y;
reg      [7:0] arg_0_TDATA;
reg            arg_0_TVALID;
reg            arg_1_TREADY;
reg    [647:0] proc_in;
reg     [71:0] stencil_0;
reg     [71:0] stencil_1;
reg     [71:0] stencil_2;
reg     [71:0] stencil_3;
reg     [71:0] stencil_4;
reg     [71:0] stencil_5;
reg     [71:0] stencil_6;
reg     [71:0] stencil_7;
reg     [71:0] stencil_8;
wire            arg_0_TREADY;
wire      [7:0] arg_1_TDATA;
wire            arg_1_TVALID;
wire            n0;
wire            n1;
wire            n2;
wire            n3;
wire      [2:0] n4;
wire      [2:0] n5;
wire      [2:0] n6;
wire      [2:0] n7;
wire      [2:0] n8;
wire      [8:0] n9;
wire      [8:0] n10;
wire      [8:0] n11;
wire      [8:0] n12;
wire            n13;
wire      [9:0] n14;
wire      [9:0] n15;
wire      [9:0] n16;
wire      [9:0] n17;
wire      [9:0] n18;
wire            n19;
wire      [7:0] n20;
wire      [7:0] n21;
wire      [7:0] n22;
wire      [7:0] n23;
wire      [7:0] n24;
wire      [7:0] n25;
wire      [7:0] n26;
wire      [7:0] n27;
wire      [7:0] n28;
wire     [15:0] n29;
wire     [23:0] n30;
wire     [31:0] n31;
wire     [39:0] n32;
wire     [47:0] n33;
wire     [55:0] n34;
wire     [63:0] n35;
wire     [71:0] n36;
wire      [7:0] n37;
wire      [7:0] n38;
wire      [7:0] n39;
wire      [7:0] n40;
wire      [7:0] n41;
wire      [7:0] n42;
wire      [7:0] n43;
wire      [7:0] n44;
wire      [7:0] n45;
wire     [15:0] n46;
wire     [23:0] n47;
wire     [31:0] n48;
wire     [39:0] n49;
wire     [47:0] n50;
wire     [55:0] n51;
wire     [63:0] n52;
wire     [71:0] n53;
wire      [7:0] n54;
wire      [7:0] n55;
wire      [7:0] n56;
wire      [7:0] n57;
wire      [7:0] n58;
wire      [7:0] n59;
wire      [7:0] n60;
wire      [7:0] n61;
wire      [7:0] n62;
wire     [15:0] n63;
wire     [23:0] n64;
wire     [31:0] n65;
wire     [39:0] n66;
wire     [47:0] n67;
wire     [55:0] n68;
wire     [63:0] n69;
wire     [71:0] n70;
wire      [7:0] n71;
wire      [7:0] n72;
wire      [7:0] n73;
wire      [7:0] n74;
wire      [7:0] n75;
wire      [7:0] n76;
wire      [7:0] n77;
wire      [7:0] n78;
wire      [7:0] n79;
wire     [15:0] n80;
wire     [23:0] n81;
wire     [31:0] n82;
wire     [39:0] n83;
wire     [47:0] n84;
wire     [55:0] n85;
wire     [63:0] n86;
wire     [71:0] n87;
wire      [7:0] n88;
wire      [7:0] n89;
wire      [7:0] n90;
wire      [7:0] n91;
wire      [7:0] n92;
wire      [7:0] n93;
wire      [7:0] n94;
wire      [7:0] n95;
wire      [7:0] n96;
wire     [15:0] n97;
wire     [23:0] n98;
wire     [31:0] n99;
wire     [39:0] n100;
wire     [47:0] n101;
wire     [55:0] n102;
wire     [63:0] n103;
wire     [71:0] n104;
wire      [7:0] n105;
wire      [7:0] n106;
wire      [7:0] n107;
wire      [7:0] n108;
wire      [7:0] n109;
wire      [7:0] n110;
wire      [7:0] n111;
wire      [7:0] n112;
wire      [7:0] n113;
wire     [15:0] n114;
wire     [23:0] n115;
wire     [31:0] n116;
wire     [39:0] n117;
wire     [47:0] n118;
wire     [55:0] n119;
wire     [63:0] n120;
wire     [71:0] n121;
wire      [7:0] n122;
wire      [7:0] n123;
wire      [7:0] n124;
wire      [7:0] n125;
wire      [7:0] n126;
wire      [7:0] n127;
wire      [7:0] n128;
wire      [7:0] n129;
wire      [7:0] n130;
wire     [15:0] n131;
wire     [23:0] n132;
wire     [31:0] n133;
wire     [39:0] n134;
wire     [47:0] n135;
wire     [55:0] n136;
wire     [63:0] n137;
wire     [71:0] n138;
wire      [7:0] n139;
wire      [7:0] n140;
wire      [7:0] n141;
wire      [7:0] n142;
wire      [7:0] n143;
wire      [7:0] n144;
wire      [7:0] n145;
wire      [7:0] n146;
wire      [7:0] n147;
wire     [15:0] n148;
wire     [23:0] n149;
wire     [31:0] n150;
wire     [39:0] n151;
wire     [47:0] n152;
wire     [55:0] n153;
wire     [63:0] n154;
wire     [71:0] n155;
wire      [7:0] n156;
wire      [7:0] n157;
wire      [7:0] n158;
wire      [7:0] n159;
wire      [7:0] n160;
wire      [7:0] n161;
wire      [7:0] n162;
wire      [7:0] n163;
wire      [7:0] n164;
wire     [15:0] n165;
wire     [23:0] n166;
wire     [31:0] n167;
wire     [39:0] n168;
wire     [47:0] n169;
wire     [55:0] n170;
wire     [63:0] n171;
wire     [71:0] n172;
wire    [143:0] n173;
wire    [215:0] n174;
wire    [287:0] n175;
wire    [359:0] n176;
wire    [431:0] n177;
wire    [503:0] n178;
wire    [575:0] n179;
wire    [647:0] n180;
wire    [647:0] n181;
wire      [7:0] n182;
wire      [7:0] n183;
wire      [7:0] n184;
wire            n185;
wire            n186;
wire            n187;
wire            n188;
wire            n189;
wire    [647:0] n190;
wire            n191;
wire     [71:0] n192;
wire     [71:0] n193;
wire     [71:0] n194;
wire     [71:0] n195;
wire     [71:0] n196;
wire     [71:0] n197;
wire     [71:0] n198;
wire     [71:0] n199;
wire     [71:0] n200;
wire     [71:0] n201;
wire     [71:0] n202;
wire     [71:0] n203;
wire     [71:0] n204;
wire     [71:0] n205;
wire     [71:0] n206;
wire     [71:0] n207;
wire     [71:0] n208;
wire     [71:0] n209;
wire     [71:0] n210;
wire     [71:0] n211;
wire     [71:0] n212;
wire     [71:0] n213;
wire     [71:0] n214;
wire     [71:0] n215;
wire            n216;
wire      [8:0] n217;
wire      [7:0] n218;
wire            n219;
wire            n220;
wire            n221;
wire            n222;
wire            n223;
wire            n224;
wire      [7:0] n225;
wire      [7:0] n226;
wire      [7:0] n227;
wire      [7:0] n228;
wire      [7:0] n229;
wire      [7:0] n230;
wire      [7:0] n231;
wire      [7:0] n232;
wire      [7:0] n233;
wire      [7:0] n234;
wire      [7:0] n235;
wire      [7:0] n236;
wire      [7:0] n237;
wire      [7:0] n238;
wire      [7:0] n239;
wire      [7:0] n240;
wire      [7:0] n241;
wire      [7:0] n242;
wire      [7:0] n243;
wire      [7:0] n244;
wire      [7:0] n245;
wire      [7:0] n246;
wire      [7:0] n247;
wire      [7:0] n248;
wire      [7:0] n249;
wire      [7:0] n250;
wire      [7:0] n251;
wire      [7:0] n252;
wire      [7:0] n253;
wire      [7:0] n254;
wire      [7:0] n255;
wire      [7:0] n256;
wire      [7:0] n257;
wire      [7:0] n258;
wire      [7:0] n259;
wire      [7:0] n260;
wire      [7:0] n261;
wire      [7:0] n262;
wire      [7:0] n263;
wire      [7:0] n264;
wire      [7:0] n265;
wire      [7:0] n266;
wire      [7:0] n267;
wire      [7:0] n268;
wire      [7:0] n269;
wire      [7:0] n270;
wire      [7:0] n271;
wire      [7:0] n272;
wire      [7:0] n273;
wire      [7:0] n274;
wire      [7:0] n275;
wire      [7:0] n276;
wire      [7:0] n277;
wire      [7:0] n278;
wire      [7:0] n279;
wire      [7:0] n280;
wire      [7:0] n281;
wire      [7:0] n282;
wire      [7:0] n283;
wire      [7:0] n284;
wire      [7:0] n285;
wire      [7:0] n286;
wire      [7:0] n287;
wire     [15:0] n288;
wire     [23:0] n289;
wire     [31:0] n290;
wire     [39:0] n291;
wire     [47:0] n292;
wire     [55:0] n293;
wire     [63:0] n294;
wire     [71:0] n295;
wire     [71:0] n296;
wire     [71:0] n297;
wire     [71:0] n298;
wire      [8:0] RAM_0_addr0;
wire      [7:0] RAM_0_data0;
wire            n299;
wire            n300;
wire            n301;
wire            n302;
wire            n303;
wire            n304;
wire      [8:0] RAM_1_addr0;
wire      [7:0] RAM_1_data0;
wire            n305;
wire            n306;
wire            n307;
wire      [8:0] RAM_2_addr0;
wire      [7:0] RAM_2_data0;
wire            n308;
wire            n309;
wire            n310;
wire      [8:0] RAM_3_addr0;
wire      [7:0] RAM_3_data0;
wire            n311;
wire            n312;
wire            n313;
wire      [8:0] RAM_4_addr0;
wire      [7:0] RAM_4_data0;
wire            n314;
wire            n315;
wire            n316;
wire      [8:0] RAM_5_addr0;
wire      [7:0] RAM_5_data0;
wire            n317;
wire            n318;
wire            n319;
wire      [8:0] RAM_6_addr0;
wire      [7:0] RAM_6_data0;
wire            n320;
wire            n321;
wire            n322;
wire      [8:0] RAM_7_addr0;
wire      [7:0] RAM_7_data0;
wire            n323;
wire            n324;
wire            n325;
reg      [7:0] RAM_0[511:0];
reg      [7:0] RAM_1[511:0];
reg      [7:0] RAM_2[511:0];
reg      [7:0] RAM_3[511:0];
reg      [7:0] RAM_4[511:0];
reg      [7:0] RAM_5[511:0];
reg      [7:0] RAM_6[511:0];
reg      [7:0] RAM_7[511:0];
wire clk;
wire rst;
wire step;
assign n0 =  ( 1'd0 ) & ( arg_0_TREADY )  ;
assign n1 =  ( n0 ) == ( 1'd0 )  ;
assign n2 =  ( RAM_x ) == ( 9'd488 )  ;
assign n3 =  ( RAM_w ) == ( 3'd7 )  ;
assign n4 =  ( RAM_w ) + ( 3'd1 )  ;
assign n5 =  ( n3 ) ? ( 3'd0 ) : ( n4 ) ;
assign n6 =  ( n2 ) ? ( n5 ) : ( RAM_w ) ;
assign n7 =  ( n1 ) ? ( n6 ) : ( RAM_w ) ;
assign n8 =  ( n1 ) ? ( RAM_w ) : ( n7 ) ;
assign n9 =  ( RAM_x ) + ( 9'd1 )  ;
assign n10 =  ( n2 ) ? ( 9'd1 ) : ( n9 ) ;
assign n11 =  ( n1 ) ? ( n10 ) : ( RAM_x ) ;
assign n12 =  ( n1 ) ? ( RAM_x ) : ( n11 ) ;
assign n13 =  ( RAM_y ) == ( 10'd648 )  ;
assign n14 =  ( RAM_y ) + ( 10'd1 )  ;
assign n15 =  ( n13 ) ? ( 10'd0 ) : ( n14 ) ;
assign n16 =  ( n2 ) ? ( n15 ) : ( RAM_y ) ;
assign n17 =  ( n1 ) ? ( n16 ) : ( RAM_y ) ;
assign n18 =  ( n1 ) ? ( RAM_y ) : ( n17 ) ;
assign n19 =  ( RAM_x ) > ( 9'd9 )  ;
assign n20 = stencil_8[71:64] ;
assign n21 = stencil_7[71:64] ;
assign n22 = stencil_6[71:64] ;
assign n23 = stencil_5[71:64] ;
assign n24 = stencil_4[71:64] ;
assign n25 = stencil_3[71:64] ;
assign n26 = stencil_2[71:64] ;
assign n27 = stencil_1[71:64] ;
assign n28 = stencil_0[71:64] ;
assign n29 =  { ( n27 ) , ( n28 ) }  ;
assign n30 =  { ( n26 ) , ( n29 ) }  ;
assign n31 =  { ( n25 ) , ( n30 ) }  ;
assign n32 =  { ( n24 ) , ( n31 ) }  ;
assign n33 =  { ( n23 ) , ( n32 ) }  ;
assign n34 =  { ( n22 ) , ( n33 ) }  ;
assign n35 =  { ( n21 ) , ( n34 ) }  ;
assign n36 =  { ( n20 ) , ( n35 ) }  ;
assign n37 = stencil_8[63:56] ;
assign n38 = stencil_7[63:56] ;
assign n39 = stencil_6[63:56] ;
assign n40 = stencil_5[63:56] ;
assign n41 = stencil_4[63:56] ;
assign n42 = stencil_3[63:56] ;
assign n43 = stencil_2[63:56] ;
assign n44 = stencil_1[63:56] ;
assign n45 = stencil_0[63:56] ;
assign n46 =  { ( n44 ) , ( n45 ) }  ;
assign n47 =  { ( n43 ) , ( n46 ) }  ;
assign n48 =  { ( n42 ) , ( n47 ) }  ;
assign n49 =  { ( n41 ) , ( n48 ) }  ;
assign n50 =  { ( n40 ) , ( n49 ) }  ;
assign n51 =  { ( n39 ) , ( n50 ) }  ;
assign n52 =  { ( n38 ) , ( n51 ) }  ;
assign n53 =  { ( n37 ) , ( n52 ) }  ;
assign n54 = stencil_8[55:48] ;
assign n55 = stencil_7[55:48] ;
assign n56 = stencil_6[55:48] ;
assign n57 = stencil_5[55:48] ;
assign n58 = stencil_4[55:48] ;
assign n59 = stencil_3[55:48] ;
assign n60 = stencil_2[55:48] ;
assign n61 = stencil_1[55:48] ;
assign n62 = stencil_0[55:48] ;
assign n63 =  { ( n61 ) , ( n62 ) }  ;
assign n64 =  { ( n60 ) , ( n63 ) }  ;
assign n65 =  { ( n59 ) , ( n64 ) }  ;
assign n66 =  { ( n58 ) , ( n65 ) }  ;
assign n67 =  { ( n57 ) , ( n66 ) }  ;
assign n68 =  { ( n56 ) , ( n67 ) }  ;
assign n69 =  { ( n55 ) , ( n68 ) }  ;
assign n70 =  { ( n54 ) , ( n69 ) }  ;
assign n71 = stencil_8[47:40] ;
assign n72 = stencil_7[47:40] ;
assign n73 = stencil_6[47:40] ;
assign n74 = stencil_5[47:40] ;
assign n75 = stencil_4[47:40] ;
assign n76 = stencil_3[47:40] ;
assign n77 = stencil_2[47:40] ;
assign n78 = stencil_1[47:40] ;
assign n79 = stencil_0[47:40] ;
assign n80 =  { ( n78 ) , ( n79 ) }  ;
assign n81 =  { ( n77 ) , ( n80 ) }  ;
assign n82 =  { ( n76 ) , ( n81 ) }  ;
assign n83 =  { ( n75 ) , ( n82 ) }  ;
assign n84 =  { ( n74 ) , ( n83 ) }  ;
assign n85 =  { ( n73 ) , ( n84 ) }  ;
assign n86 =  { ( n72 ) , ( n85 ) }  ;
assign n87 =  { ( n71 ) , ( n86 ) }  ;
assign n88 = stencil_8[39:32] ;
assign n89 = stencil_7[39:32] ;
assign n90 = stencil_6[39:32] ;
assign n91 = stencil_5[39:32] ;
assign n92 = stencil_4[39:32] ;
assign n93 = stencil_3[39:32] ;
assign n94 = stencil_2[39:32] ;
assign n95 = stencil_1[39:32] ;
assign n96 = stencil_0[39:32] ;
assign n97 =  { ( n95 ) , ( n96 ) }  ;
assign n98 =  { ( n94 ) , ( n97 ) }  ;
assign n99 =  { ( n93 ) , ( n98 ) }  ;
assign n100 =  { ( n92 ) , ( n99 ) }  ;
assign n101 =  { ( n91 ) , ( n100 ) }  ;
assign n102 =  { ( n90 ) , ( n101 ) }  ;
assign n103 =  { ( n89 ) , ( n102 ) }  ;
assign n104 =  { ( n88 ) , ( n103 ) }  ;
assign n105 = stencil_8[31:24] ;
assign n106 = stencil_7[31:24] ;
assign n107 = stencil_6[31:24] ;
assign n108 = stencil_5[31:24] ;
assign n109 = stencil_4[31:24] ;
assign n110 = stencil_3[31:24] ;
assign n111 = stencil_2[31:24] ;
assign n112 = stencil_1[31:24] ;
assign n113 = stencil_0[31:24] ;
assign n114 =  { ( n112 ) , ( n113 ) }  ;
assign n115 =  { ( n111 ) , ( n114 ) }  ;
assign n116 =  { ( n110 ) , ( n115 ) }  ;
assign n117 =  { ( n109 ) , ( n116 ) }  ;
assign n118 =  { ( n108 ) , ( n117 ) }  ;
assign n119 =  { ( n107 ) , ( n118 ) }  ;
assign n120 =  { ( n106 ) , ( n119 ) }  ;
assign n121 =  { ( n105 ) , ( n120 ) }  ;
assign n122 = stencil_8[23:16] ;
assign n123 = stencil_7[23:16] ;
assign n124 = stencil_6[23:16] ;
assign n125 = stencil_5[23:16] ;
assign n126 = stencil_4[23:16] ;
assign n127 = stencil_3[23:16] ;
assign n128 = stencil_2[23:16] ;
assign n129 = stencil_1[23:16] ;
assign n130 = stencil_0[23:16] ;
assign n131 =  { ( n129 ) , ( n130 ) }  ;
assign n132 =  { ( n128 ) , ( n131 ) }  ;
assign n133 =  { ( n127 ) , ( n132 ) }  ;
assign n134 =  { ( n126 ) , ( n133 ) }  ;
assign n135 =  { ( n125 ) , ( n134 ) }  ;
assign n136 =  { ( n124 ) , ( n135 ) }  ;
assign n137 =  { ( n123 ) , ( n136 ) }  ;
assign n138 =  { ( n122 ) , ( n137 ) }  ;
assign n139 = stencil_8[15:8] ;
assign n140 = stencil_7[15:8] ;
assign n141 = stencil_6[15:8] ;
assign n142 = stencil_5[15:8] ;
assign n143 = stencil_4[15:8] ;
assign n144 = stencil_3[15:8] ;
assign n145 = stencil_2[15:8] ;
assign n146 = stencil_1[15:8] ;
assign n147 = stencil_0[15:8] ;
assign n148 =  { ( n146 ) , ( n147 ) }  ;
assign n149 =  { ( n145 ) , ( n148 ) }  ;
assign n150 =  { ( n144 ) , ( n149 ) }  ;
assign n151 =  { ( n143 ) , ( n150 ) }  ;
assign n152 =  { ( n142 ) , ( n151 ) }  ;
assign n153 =  { ( n141 ) , ( n152 ) }  ;
assign n154 =  { ( n140 ) , ( n153 ) }  ;
assign n155 =  { ( n139 ) , ( n154 ) }  ;
assign n156 = stencil_8[7:0] ;
assign n157 = stencil_7[7:0] ;
assign n158 = stencil_6[7:0] ;
assign n159 = stencil_5[7:0] ;
assign n160 = stencil_4[7:0] ;
assign n161 = stencil_3[7:0] ;
assign n162 = stencil_2[7:0] ;
assign n163 = stencil_1[7:0] ;
assign n164 = stencil_0[7:0] ;
assign n165 =  { ( n163 ) , ( n164 ) }  ;
assign n166 =  { ( n162 ) , ( n165 ) }  ;
assign n167 =  { ( n161 ) , ( n166 ) }  ;
assign n168 =  { ( n160 ) , ( n167 ) }  ;
assign n169 =  { ( n159 ) , ( n168 ) }  ;
assign n170 =  { ( n158 ) , ( n169 ) }  ;
assign n171 =  { ( n157 ) , ( n170 ) }  ;
assign n172 =  { ( n156 ) , ( n171 ) }  ;
assign n173 =  { ( n155 ) , ( n172 ) }  ;
assign n174 =  { ( n138 ) , ( n173 ) }  ;
assign n175 =  { ( n121 ) , ( n174 ) }  ;
assign n176 =  { ( n104 ) , ( n175 ) }  ;
assign n177 =  { ( n87 ) , ( n176 ) }  ;
assign n178 =  { ( n70 ) , ( n177 ) }  ;
assign n179 =  { ( n53 ) , ( n178 ) }  ;
assign n180 =  { ( n36 ) , ( n179 ) }  ;
assign n181 =  ( n19 ) ? ( n180 ) : ( proc_in ) ;
assign n182 = gb_fun(n181) ;
assign n183 =  ( n1 ) ? ( arg_0_TDATA ) : ( arg_0_TDATA ) ;
assign n184 =  ( n1 ) ? ( n182 ) : ( n183 ) ;
assign n185 =  ( n19 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n186 =  ( n1 ) ? ( 1'd0 ) : ( arg_0_TVALID ) ;
assign n187 =  ( n1 ) ? ( n185 ) : ( n186 ) ;
assign n188 =  ( n1 ) ? ( 1'd0 ) : ( arg_1_TREADY ) ;
assign n189 =  ( n1 ) ? ( 1'd1 ) : ( n188 ) ;
assign n190 =  ( n1 ) ? ( n181 ) : ( proc_in ) ;
assign n191 =  ( RAM_y ) < ( 10'd8 )  ;
assign n192 =  ( n191 ) ? ( stencil_0 ) : ( stencil_1 ) ;
assign n193 =  ( n1 ) ? ( stencil_0 ) : ( stencil_0 ) ;
assign n194 =  ( n1 ) ? ( n192 ) : ( n193 ) ;
assign n195 =  ( n191 ) ? ( stencil_1 ) : ( stencil_2 ) ;
assign n196 =  ( n1 ) ? ( stencil_1 ) : ( stencil_1 ) ;
assign n197 =  ( n1 ) ? ( n195 ) : ( n196 ) ;
assign n198 =  ( n191 ) ? ( stencil_2 ) : ( stencil_3 ) ;
assign n199 =  ( n1 ) ? ( stencil_2 ) : ( stencil_2 ) ;
assign n200 =  ( n1 ) ? ( n198 ) : ( n199 ) ;
assign n201 =  ( n191 ) ? ( stencil_3 ) : ( stencil_4 ) ;
assign n202 =  ( n1 ) ? ( stencil_3 ) : ( stencil_3 ) ;
assign n203 =  ( n1 ) ? ( n201 ) : ( n202 ) ;
assign n204 =  ( n191 ) ? ( stencil_4 ) : ( stencil_5 ) ;
assign n205 =  ( n1 ) ? ( stencil_4 ) : ( stencil_4 ) ;
assign n206 =  ( n1 ) ? ( n204 ) : ( n205 ) ;
assign n207 =  ( n191 ) ? ( stencil_5 ) : ( stencil_6 ) ;
assign n208 =  ( n1 ) ? ( stencil_5 ) : ( stencil_5 ) ;
assign n209 =  ( n1 ) ? ( n207 ) : ( n208 ) ;
assign n210 =  ( n191 ) ? ( stencil_6 ) : ( stencil_7 ) ;
assign n211 =  ( n1 ) ? ( stencil_6 ) : ( stencil_6 ) ;
assign n212 =  ( n1 ) ? ( n210 ) : ( n211 ) ;
assign n213 =  ( n191 ) ? ( stencil_7 ) : ( stencil_8 ) ;
assign n214 =  ( n1 ) ? ( stencil_7 ) : ( stencil_7 ) ;
assign n215 =  ( n1 ) ? ( n213 ) : ( n214 ) ;
assign n216 =  ( RAM_w ) == ( 3'd0 )  ;
assign n217 =  ( RAM_x ) - ( 9'd1 )  ;
assign n218 =  (  RAM_7 [ n217 ] )  ;
assign n219 =  ( RAM_w ) == ( 3'd1 )  ;
assign n220 =  ( RAM_w ) == ( 3'd2 )  ;
assign n221 =  ( RAM_w ) == ( 3'd3 )  ;
assign n222 =  ( RAM_w ) == ( 3'd4 )  ;
assign n223 =  ( RAM_w ) == ( 3'd5 )  ;
assign n224 =  ( RAM_w ) == ( 3'd6 )  ;
assign n225 =  (  RAM_6 [ n217 ] )  ;
assign n226 =  ( n224 ) ? ( n218 ) : ( n225 ) ;
assign n227 =  ( n223 ) ? ( n218 ) : ( n226 ) ;
assign n228 =  ( n222 ) ? ( n218 ) : ( n227 ) ;
assign n229 =  ( n221 ) ? ( n218 ) : ( n228 ) ;
assign n230 =  ( n220 ) ? ( n218 ) : ( n229 ) ;
assign n231 =  ( n219 ) ? ( n218 ) : ( n230 ) ;
assign n232 =  ( n216 ) ? ( n218 ) : ( n231 ) ;
assign n233 =  (  RAM_5 [ n217 ] )  ;
assign n234 =  ( n224 ) ? ( n225 ) : ( n233 ) ;
assign n235 =  ( n223 ) ? ( n225 ) : ( n234 ) ;
assign n236 =  ( n222 ) ? ( n225 ) : ( n235 ) ;
assign n237 =  ( n221 ) ? ( n225 ) : ( n236 ) ;
assign n238 =  ( n220 ) ? ( n225 ) : ( n237 ) ;
assign n239 =  ( n219 ) ? ( n225 ) : ( n238 ) ;
assign n240 =  ( n216 ) ? ( n225 ) : ( n239 ) ;
assign n241 =  (  RAM_4 [ n217 ] )  ;
assign n242 =  ( n224 ) ? ( n233 ) : ( n241 ) ;
assign n243 =  ( n223 ) ? ( n233 ) : ( n242 ) ;
assign n244 =  ( n222 ) ? ( n233 ) : ( n243 ) ;
assign n245 =  ( n221 ) ? ( n233 ) : ( n244 ) ;
assign n246 =  ( n220 ) ? ( n233 ) : ( n245 ) ;
assign n247 =  ( n219 ) ? ( n233 ) : ( n246 ) ;
assign n248 =  ( n216 ) ? ( n233 ) : ( n247 ) ;
assign n249 =  (  RAM_3 [ n217 ] )  ;
assign n250 =  ( n224 ) ? ( n241 ) : ( n249 ) ;
assign n251 =  ( n223 ) ? ( n241 ) : ( n250 ) ;
assign n252 =  ( n222 ) ? ( n241 ) : ( n251 ) ;
assign n253 =  ( n221 ) ? ( n241 ) : ( n252 ) ;
assign n254 =  ( n220 ) ? ( n241 ) : ( n253 ) ;
assign n255 =  ( n219 ) ? ( n241 ) : ( n254 ) ;
assign n256 =  ( n216 ) ? ( n241 ) : ( n255 ) ;
assign n257 =  (  RAM_2 [ n217 ] )  ;
assign n258 =  ( n224 ) ? ( n249 ) : ( n257 ) ;
assign n259 =  ( n223 ) ? ( n249 ) : ( n258 ) ;
assign n260 =  ( n222 ) ? ( n249 ) : ( n259 ) ;
assign n261 =  ( n221 ) ? ( n249 ) : ( n260 ) ;
assign n262 =  ( n220 ) ? ( n249 ) : ( n261 ) ;
assign n263 =  ( n219 ) ? ( n249 ) : ( n262 ) ;
assign n264 =  ( n216 ) ? ( n249 ) : ( n263 ) ;
assign n265 =  (  RAM_1 [ n217 ] )  ;
assign n266 =  ( n224 ) ? ( n257 ) : ( n265 ) ;
assign n267 =  ( n223 ) ? ( n257 ) : ( n266 ) ;
assign n268 =  ( n222 ) ? ( n257 ) : ( n267 ) ;
assign n269 =  ( n221 ) ? ( n257 ) : ( n268 ) ;
assign n270 =  ( n220 ) ? ( n257 ) : ( n269 ) ;
assign n271 =  ( n219 ) ? ( n257 ) : ( n270 ) ;
assign n272 =  ( n216 ) ? ( n257 ) : ( n271 ) ;
assign n273 =  (  RAM_0 [ n217 ] )  ;
assign n274 =  ( n224 ) ? ( n265 ) : ( n273 ) ;
assign n275 =  ( n223 ) ? ( n265 ) : ( n274 ) ;
assign n276 =  ( n222 ) ? ( n265 ) : ( n275 ) ;
assign n277 =  ( n221 ) ? ( n265 ) : ( n276 ) ;
assign n278 =  ( n220 ) ? ( n265 ) : ( n277 ) ;
assign n279 =  ( n219 ) ? ( n265 ) : ( n278 ) ;
assign n280 =  ( n216 ) ? ( n265 ) : ( n279 ) ;
assign n281 =  ( n224 ) ? ( n273 ) : ( n218 ) ;
assign n282 =  ( n223 ) ? ( n273 ) : ( n281 ) ;
assign n283 =  ( n222 ) ? ( n273 ) : ( n282 ) ;
assign n284 =  ( n221 ) ? ( n273 ) : ( n283 ) ;
assign n285 =  ( n220 ) ? ( n273 ) : ( n284 ) ;
assign n286 =  ( n219 ) ? ( n273 ) : ( n285 ) ;
assign n287 =  ( n216 ) ? ( n273 ) : ( n286 ) ;
assign n288 =  { ( n280 ) , ( n287 ) }  ;
assign n289 =  { ( n272 ) , ( n288 ) }  ;
assign n290 =  { ( n264 ) , ( n289 ) }  ;
assign n291 =  { ( n256 ) , ( n290 ) }  ;
assign n292 =  { ( n248 ) , ( n291 ) }  ;
assign n293 =  { ( n240 ) , ( n292 ) }  ;
assign n294 =  { ( n232 ) , ( n293 ) }  ;
assign n295 =  { ( arg_1_TDATA ) , ( n294 ) }  ;
assign n296 =  ( n191 ) ? ( stencil_8 ) : ( n295 ) ;
assign n297 =  ( n1 ) ? ( n296 ) : ( stencil_8 ) ;
assign n298 =  ( n1 ) ? ( stencil_8 ) : ( n297 ) ;
assign n299 = ~ ( n1 ) ;
assign n300 =  ( n299 ) & ( n299 )  ;
assign n301 =  ( n299 ) & ( n1 )  ;
assign n302 = ~ ( n216 ) ;
assign n303 =  ( n301 ) & ( n302 )  ;
assign n304 =  ( n301 ) & ( n216 )  ;
assign RAM_0_addr0 = n304 ? (n217) : (0);
assign RAM_0_data0 = n304 ? (arg_1_TDATA) : (RAM_0[0]);
assign n305 = ~ ( n219 ) ;
assign n306 =  ( n301 ) & ( n305 )  ;
assign n307 =  ( n301 ) & ( n219 )  ;
assign RAM_1_addr0 = n307 ? (n217) : (0);
assign RAM_1_data0 = n307 ? (arg_1_TDATA) : (RAM_1[0]);
assign n308 = ~ ( n220 ) ;
assign n309 =  ( n301 ) & ( n308 )  ;
assign n310 =  ( n301 ) & ( n220 )  ;
assign RAM_2_addr0 = n310 ? (n217) : (0);
assign RAM_2_data0 = n310 ? (arg_1_TDATA) : (RAM_2[0]);
assign n311 = ~ ( n221 ) ;
assign n312 =  ( n301 ) & ( n311 )  ;
assign n313 =  ( n301 ) & ( n221 )  ;
assign RAM_3_addr0 = n313 ? (n217) : (0);
assign RAM_3_data0 = n313 ? (arg_1_TDATA) : (RAM_3[0]);
assign n314 = ~ ( n222 ) ;
assign n315 =  ( n301 ) & ( n314 )  ;
assign n316 =  ( n301 ) & ( n222 )  ;
assign RAM_4_addr0 = n316 ? (n217) : (0);
assign RAM_4_data0 = n316 ? (arg_1_TDATA) : (RAM_4[0]);
assign n317 = ~ ( n223 ) ;
assign n318 =  ( n301 ) & ( n317 )  ;
assign n319 =  ( n301 ) & ( n223 )  ;
assign RAM_5_addr0 = n319 ? (n217) : (0);
assign RAM_5_data0 = n319 ? (arg_1_TDATA) : (RAM_5[0]);
assign n320 = ~ ( n224 ) ;
assign n321 =  ( n301 ) & ( n320 )  ;
assign n322 =  ( n301 ) & ( n224 )  ;
assign RAM_6_addr0 = n322 ? (n217) : (0);
assign RAM_6_data0 = n322 ? (arg_1_TDATA) : (RAM_6[0]);
assign n323 = ~ ( n3 ) ;
assign n324 =  ( n301 ) & ( n323 )  ;
assign n325 =  ( n301 ) & ( n3 )  ;
assign RAM_7_addr0 = n325 ? (n217) : (0);
assign RAM_7_data0 = n325 ? (arg_1_TDATA) : (RAM_7[0]);
function [7:0] gb_fun ;
input [647:0] arg0;
    begin
//TODO: Add the specific function HERE.    end
endfunction

always @(posedge clk) begin
   if(rst) begin
       RAM_w <= RAM_w;
       RAM_x <= RAM_x;
       RAM_y <= RAM_y;
       arg_0_TDATA <= arg_0_TDATA;
       arg_0_TVALID <= arg_0_TVALID;
       arg_1_TREADY <= arg_1_TREADY;
       proc_in <= proc_in;
       stencil_0 <= stencil_0;
       stencil_1 <= stencil_1;
       stencil_2 <= stencil_2;
       stencil_3 <= stencil_3;
       stencil_4 <= stencil_4;
       stencil_5 <= stencil_5;
       stencil_6 <= stencil_6;
       stencil_7 <= stencil_7;
       stencil_8 <= stencil_8;
   end
   else if(step) begin
       RAM_w <= n8;
       RAM_x <= n12;
       RAM_y <= n18;
       arg_0_TDATA <= n184;
       arg_0_TVALID <= n187;
       arg_1_TREADY <= n189;
       proc_in <= n190;
       stencil_0 <= n194;
       stencil_1 <= n197;
       stencil_2 <= n200;
       stencil_3 <= n203;
       stencil_4 <= n206;
       stencil_5 <= n209;
       stencil_6 <= n212;
       stencil_7 <= n215;
       stencil_8 <= n298;
       RAM_0 [ RAM_0_addr0 ] <= RAM_0_data0;
       RAM_1 [ RAM_1_addr0 ] <= RAM_1_data0;
       RAM_2 [ RAM_2_addr0 ] <= RAM_2_data0;
       RAM_3 [ RAM_3_addr0 ] <= RAM_3_data0;
       RAM_4 [ RAM_4_addr0 ] <= RAM_4_data0;
       RAM_5 [ RAM_5_addr0 ] <= RAM_5_data0;
       RAM_6 [ RAM_6_addr0 ] <= RAM_6_data0;
       RAM_7 [ RAM_7_addr0 ] <= RAM_7_data0;
   end
end
endmodule
