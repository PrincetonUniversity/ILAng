module SPEC_B(
arg_0_TREADY,
arg_1_TDATA,
arg_1_TVALID,
LB1D_buff,
LB1D_in,
LB1D_it_1,
LB1D_p_cnt,
LB1D_uIn,
LB2D_proc_w,
LB2D_proc_x,
LB2D_proc_y,
LB2D_shift_0,
LB2D_shift_1,
LB2D_shift_2,
LB2D_shift_3,
LB2D_shift_4,
LB2D_shift_5,
LB2D_shift_6,
LB2D_shift_7,
LB2D_shift_x,
LB2D_shift_y,
arg_0_TDATA,
arg_0_TVALID,
arg_1_TREADY,
gb_exit_it_1,
gb_exit_it_2,
gb_exit_it_3,
gb_exit_it_4,
gb_exit_it_5,
gb_exit_it_6,
gb_exit_it_7,
gb_exit_it_8,
gb_p_cnt,
gb_pp_it_1,
gb_pp_it_2,
gb_pp_it_3,
gb_pp_it_4,
gb_pp_it_5,
gb_pp_it_6,
gb_pp_it_7,
gb_pp_it_8,
gb_pp_it_9,
in_stream_buff_0,
in_stream_buff_1,
in_stream_empty,
in_stream_full,
slice_stream_buff_0,
slice_stream_buff_1,
slice_stream_empty,
slice_stream_full,
stencil_stream_buff_0,
stencil_stream_buff_1,
stencil_stream_empty,
stencil_stream_full,
clk,rst,
step
);
input            arg_0_TREADY;
input      [7:0] arg_1_TDATA;
input            arg_1_TVALID;
input clk;
input rst;
input step;
output      [7:0] LB1D_buff;
output      [7:0] LB1D_in;
output            LB1D_it_1;
output     [18:0] LB1D_p_cnt;
output      [7:0] LB1D_uIn;
output     [63:0] LB2D_proc_w;
output      [8:0] LB2D_proc_x;
output      [9:0] LB2D_proc_y;
output     [71:0] LB2D_shift_0;
output     [71:0] LB2D_shift_1;
output     [71:0] LB2D_shift_2;
output     [71:0] LB2D_shift_3;
output     [71:0] LB2D_shift_4;
output     [71:0] LB2D_shift_5;
output     [71:0] LB2D_shift_6;
output     [71:0] LB2D_shift_7;
output      [8:0] LB2D_shift_x;
output      [9:0] LB2D_shift_y;
output      [7:0] arg_0_TDATA;
output            arg_0_TVALID;
output            arg_1_TREADY;
output            gb_exit_it_1;
output            gb_exit_it_2;
output            gb_exit_it_3;
output            gb_exit_it_4;
output            gb_exit_it_5;
output            gb_exit_it_6;
output            gb_exit_it_7;
output            gb_exit_it_8;
output     [18:0] gb_p_cnt;
output            gb_pp_it_1;
output            gb_pp_it_2;
output            gb_pp_it_3;
output            gb_pp_it_4;
output            gb_pp_it_5;
output            gb_pp_it_6;
output            gb_pp_it_7;
output            gb_pp_it_8;
output            gb_pp_it_9;
output      [7:0] in_stream_buff_0;
output      [7:0] in_stream_buff_1;
output            in_stream_empty;
output            in_stream_full;
output     [71:0] slice_stream_buff_0;
output     [71:0] slice_stream_buff_1;
output            slice_stream_empty;
output            slice_stream_full;
output    [647:0] stencil_stream_buff_0;
output    [647:0] stencil_stream_buff_1;
output            stencil_stream_empty;
output            stencil_stream_full;
reg      [7:0] LB1D_buff;
reg      [7:0] LB1D_in;
reg            LB1D_it_1;
reg     [18:0] LB1D_p_cnt;
reg      [7:0] LB1D_uIn;
reg     [63:0] LB2D_proc_w;
reg      [8:0] LB2D_proc_x;
reg      [9:0] LB2D_proc_y;
reg     [71:0] LB2D_shift_0;
reg     [71:0] LB2D_shift_1;
reg     [71:0] LB2D_shift_2;
reg     [71:0] LB2D_shift_3;
reg     [71:0] LB2D_shift_4;
reg     [71:0] LB2D_shift_5;
reg     [71:0] LB2D_shift_6;
reg     [71:0] LB2D_shift_7;
reg      [8:0] LB2D_shift_x;
reg      [9:0] LB2D_shift_y;
reg      [7:0] arg_0_TDATA;
reg            arg_0_TVALID;
reg            arg_1_TREADY;
reg            gb_exit_it_1;
reg            gb_exit_it_2;
reg            gb_exit_it_3;
reg            gb_exit_it_4;
reg            gb_exit_it_5;
reg            gb_exit_it_6;
reg            gb_exit_it_7;
reg            gb_exit_it_8;
reg     [18:0] gb_p_cnt;
reg            gb_pp_it_1;
reg            gb_pp_it_2;
reg            gb_pp_it_3;
reg            gb_pp_it_4;
reg            gb_pp_it_5;
reg            gb_pp_it_6;
reg            gb_pp_it_7;
reg            gb_pp_it_8;
reg            gb_pp_it_9;
reg      [7:0] in_stream_buff_0;
reg      [7:0] in_stream_buff_1;
reg            in_stream_empty;
reg            in_stream_full;
reg     [71:0] slice_stream_buff_0;
reg     [71:0] slice_stream_buff_1;
reg            slice_stream_empty;
reg            slice_stream_full;
reg    [647:0] stencil_stream_buff_0;
reg    [647:0] stencil_stream_buff_1;
reg            stencil_stream_empty;
reg            stencil_stream_full;
wire            arg_0_TREADY;
wire      [7:0] arg_1_TDATA;
wire            arg_1_TVALID;
wire            n0;
wire            n1;
wire            n2;
wire            n3;
wire            n4;
wire            n5;
wire            n6;
wire            n7;
wire            n8;
wire            n9;
wire            n10;
wire            n11;
wire            n12;
wire            n13;
wire            n14;
wire            n15;
wire            n16;
wire            n17;
wire            n18;
wire            n19;
wire            n20;
wire            n21;
wire            n22;
wire            n23;
wire            n24;
wire            n25;
wire            n26;
wire            n27;
wire            n28;
wire            n29;
wire            n30;
wire            n31;
wire            n32;
wire      [7:0] n33;
wire      [7:0] n34;
wire      [7:0] n35;
wire      [7:0] n36;
wire      [7:0] n37;
wire      [7:0] n38;
wire      [7:0] n39;
wire      [7:0] n40;
wire      [7:0] n41;
wire      [7:0] n42;
wire      [7:0] n43;
wire      [7:0] n44;
wire            n45;
wire     [18:0] n46;
wire     [18:0] n47;
wire            n48;
wire     [18:0] n49;
wire     [18:0] n50;
wire     [18:0] n51;
wire     [18:0] n52;
wire     [18:0] n53;
wire     [18:0] n54;
wire     [18:0] n55;
wire      [7:0] n56;
wire      [7:0] n57;
wire      [7:0] n58;
wire      [7:0] n59;
wire      [7:0] n60;
wire            n61;
wire            n62;
wire     [63:0] n63;
wire     [63:0] n64;
wire     [63:0] n65;
wire     [63:0] n66;
wire     [63:0] n67;
wire     [63:0] n68;
wire     [63:0] n69;
wire     [63:0] n70;
wire      [8:0] n71;
wire      [8:0] n72;
wire      [8:0] n73;
wire      [8:0] n74;
wire      [8:0] n75;
wire      [8:0] n76;
wire      [8:0] n77;
wire            n78;
wire      [9:0] n79;
wire      [9:0] n80;
wire      [9:0] n81;
wire      [9:0] n82;
wire      [9:0] n83;
wire      [9:0] n84;
wire      [9:0] n85;
wire      [9:0] n86;
wire     [71:0] n87;
wire     [71:0] n88;
wire     [71:0] n89;
wire     [71:0] n90;
wire     [71:0] n91;
wire     [71:0] n92;
wire     [71:0] n93;
wire     [71:0] n94;
wire     [71:0] n95;
wire     [71:0] n96;
wire     [71:0] n97;
wire     [71:0] n98;
wire     [71:0] n99;
wire     [71:0] n100;
wire     [71:0] n101;
wire     [71:0] n102;
wire     [71:0] n103;
wire     [71:0] n104;
wire     [71:0] n105;
wire     [71:0] n106;
wire     [71:0] n107;
wire     [71:0] n108;
wire     [71:0] n109;
wire     [71:0] n110;
wire     [71:0] n111;
wire     [71:0] n112;
wire     [71:0] n113;
wire     [71:0] n114;
wire     [71:0] n115;
wire     [71:0] n116;
wire     [71:0] n117;
wire     [71:0] n118;
wire     [71:0] n119;
wire     [71:0] n120;
wire     [71:0] n121;
wire            n122;
wire     [71:0] n123;
wire     [71:0] n124;
wire     [71:0] n125;
wire     [71:0] n126;
wire     [71:0] n127;
wire     [71:0] n128;
wire      [8:0] n129;
wire      [8:0] n130;
wire      [8:0] n131;
wire      [8:0] n132;
wire      [8:0] n133;
wire      [8:0] n134;
wire            n135;
wire            n136;
wire      [9:0] n137;
wire      [9:0] n138;
wire      [9:0] n139;
wire      [9:0] n140;
wire      [9:0] n141;
wire      [9:0] n142;
wire      [9:0] n143;
wire      [9:0] n144;
wire            n145;
wire    [647:0] n146;
wire      [7:0] n147;
wire      [7:0] n148;
wire      [7:0] n149;
wire      [7:0] n150;
wire      [7:0] n151;
wire      [7:0] n152;
wire            n153;
wire            n154;
wire            n155;
wire            n156;
wire            n157;
wire            n158;
wire            n159;
wire            n160;
wire            n161;
wire            n162;
wire            n163;
wire            n164;
wire            n165;
wire     [18:0] n166;
wire            n167;
wire            n168;
wire            n169;
wire            n170;
wire            n171;
wire            n172;
wire            n173;
wire            n174;
wire            n175;
wire            n176;
wire            n177;
wire            n178;
wire            n179;
wire            n180;
wire            n181;
wire            n182;
wire            n183;
wire            n184;
wire            n185;
wire            n186;
wire            n187;
wire            n188;
wire            n189;
wire            n190;
wire            n191;
wire            n192;
wire            n193;
wire            n194;
wire            n195;
wire            n196;
wire            n197;
wire            n198;
wire            n199;
wire            n200;
wire            n201;
wire            n202;
wire            n203;
wire            n204;
wire            n205;
wire            n206;
wire            n207;
wire            n208;
wire            n209;
wire     [18:0] n210;
wire     [18:0] n211;
wire     [18:0] n212;
wire     [18:0] n213;
wire     [18:0] n214;
wire     [18:0] n215;
wire            n216;
wire            n217;
wire            n218;
wire            n219;
wire            n220;
wire            n221;
wire            n222;
wire            n223;
wire            n224;
wire            n225;
wire            n226;
wire            n227;
wire            n228;
wire            n229;
wire            n230;
wire            n231;
wire            n232;
wire            n233;
wire            n234;
wire            n235;
wire            n236;
wire            n237;
wire            n238;
wire            n239;
wire            n240;
wire            n241;
wire            n242;
wire            n243;
wire            n244;
wire            n245;
wire            n246;
wire            n247;
wire            n248;
wire            n249;
wire            n250;
wire            n251;
wire            n252;
wire            n253;
wire            n254;
wire            n255;
wire            n256;
wire            n257;
wire            n258;
wire            n259;
wire            n260;
wire      [7:0] n261;
wire      [7:0] n262;
wire      [7:0] n263;
wire      [7:0] n264;
wire      [7:0] n265;
wire      [7:0] n266;
wire      [7:0] n267;
wire      [7:0] n268;
wire      [7:0] n269;
wire      [7:0] n270;
wire            n271;
wire            n272;
wire            n273;
wire            n274;
wire            n275;
wire            n276;
wire            n277;
wire            n278;
wire            n279;
wire            n280;
wire            n281;
wire            n282;
wire            n283;
wire            n284;
wire      [7:0] n285;
wire            n286;
wire      [8:0] n287;
wire      [7:0] n288;
wire            n289;
wire      [7:0] n290;
wire            n291;
wire      [7:0] n292;
wire            n293;
wire      [7:0] n294;
wire            n295;
wire      [7:0] n296;
wire            n297;
wire      [7:0] n298;
wire            n299;
wire      [7:0] n300;
wire      [7:0] n301;
wire      [7:0] n302;
wire      [7:0] n303;
wire      [7:0] n304;
wire      [7:0] n305;
wire      [7:0] n306;
wire      [7:0] n307;
wire      [7:0] n308;
wire      [7:0] n309;
wire      [7:0] n310;
wire      [7:0] n311;
wire      [7:0] n312;
wire      [7:0] n313;
wire      [7:0] n314;
wire      [7:0] n315;
wire      [7:0] n316;
wire      [7:0] n317;
wire      [7:0] n318;
wire      [7:0] n319;
wire      [7:0] n320;
wire      [7:0] n321;
wire      [7:0] n322;
wire      [7:0] n323;
wire      [7:0] n324;
wire      [7:0] n325;
wire      [7:0] n326;
wire      [7:0] n327;
wire      [7:0] n328;
wire      [7:0] n329;
wire      [7:0] n330;
wire      [7:0] n331;
wire      [7:0] n332;
wire      [7:0] n333;
wire      [7:0] n334;
wire      [7:0] n335;
wire      [7:0] n336;
wire      [7:0] n337;
wire      [7:0] n338;
wire      [7:0] n339;
wire      [7:0] n340;
wire      [7:0] n341;
wire      [7:0] n342;
wire      [7:0] n343;
wire      [7:0] n344;
wire      [7:0] n345;
wire      [7:0] n346;
wire      [7:0] n347;
wire      [7:0] n348;
wire      [7:0] n349;
wire      [7:0] n350;
wire      [7:0] n351;
wire      [7:0] n352;
wire      [7:0] n353;
wire      [7:0] n354;
wire      [7:0] n355;
wire      [7:0] n356;
wire      [7:0] n357;
wire     [15:0] n358;
wire     [23:0] n359;
wire     [31:0] n360;
wire     [39:0] n361;
wire     [47:0] n362;
wire     [55:0] n363;
wire     [63:0] n364;
wire     [71:0] n365;
wire     [71:0] n366;
wire     [71:0] n367;
wire     [71:0] n368;
wire     [71:0] n369;
wire     [71:0] n370;
wire     [71:0] n371;
wire     [71:0] n372;
wire     [71:0] n373;
wire     [71:0] n374;
wire     [71:0] n375;
wire     [71:0] n376;
wire     [71:0] n377;
wire            n378;
wire            n379;
wire            n380;
wire            n381;
wire            n382;
wire            n383;
wire            n384;
wire            n385;
wire            n386;
wire            n387;
wire            n388;
wire            n389;
wire            n390;
wire            n391;
wire            n392;
wire            n393;
wire      [7:0] n394;
wire      [7:0] n395;
wire      [7:0] n396;
wire      [7:0] n397;
wire      [7:0] n398;
wire      [7:0] n399;
wire      [7:0] n400;
wire      [7:0] n401;
wire      [7:0] n402;
wire     [15:0] n403;
wire     [23:0] n404;
wire     [31:0] n405;
wire     [39:0] n406;
wire     [47:0] n407;
wire     [55:0] n408;
wire     [63:0] n409;
wire     [71:0] n410;
wire      [7:0] n411;
wire      [7:0] n412;
wire      [7:0] n413;
wire      [7:0] n414;
wire      [7:0] n415;
wire      [7:0] n416;
wire      [7:0] n417;
wire      [7:0] n418;
wire      [7:0] n419;
wire     [15:0] n420;
wire     [23:0] n421;
wire     [31:0] n422;
wire     [39:0] n423;
wire     [47:0] n424;
wire     [55:0] n425;
wire     [63:0] n426;
wire     [71:0] n427;
wire      [7:0] n428;
wire      [7:0] n429;
wire      [7:0] n430;
wire      [7:0] n431;
wire      [7:0] n432;
wire      [7:0] n433;
wire      [7:0] n434;
wire      [7:0] n435;
wire      [7:0] n436;
wire     [15:0] n437;
wire     [23:0] n438;
wire     [31:0] n439;
wire     [39:0] n440;
wire     [47:0] n441;
wire     [55:0] n442;
wire     [63:0] n443;
wire     [71:0] n444;
wire      [7:0] n445;
wire      [7:0] n446;
wire      [7:0] n447;
wire      [7:0] n448;
wire      [7:0] n449;
wire      [7:0] n450;
wire      [7:0] n451;
wire      [7:0] n452;
wire      [7:0] n453;
wire     [15:0] n454;
wire     [23:0] n455;
wire     [31:0] n456;
wire     [39:0] n457;
wire     [47:0] n458;
wire     [55:0] n459;
wire     [63:0] n460;
wire     [71:0] n461;
wire      [7:0] n462;
wire      [7:0] n463;
wire      [7:0] n464;
wire      [7:0] n465;
wire      [7:0] n466;
wire      [7:0] n467;
wire      [7:0] n468;
wire      [7:0] n469;
wire      [7:0] n470;
wire     [15:0] n471;
wire     [23:0] n472;
wire     [31:0] n473;
wire     [39:0] n474;
wire     [47:0] n475;
wire     [55:0] n476;
wire     [63:0] n477;
wire     [71:0] n478;
wire      [7:0] n479;
wire      [7:0] n480;
wire      [7:0] n481;
wire      [7:0] n482;
wire      [7:0] n483;
wire      [7:0] n484;
wire      [7:0] n485;
wire      [7:0] n486;
wire      [7:0] n487;
wire     [15:0] n488;
wire     [23:0] n489;
wire     [31:0] n490;
wire     [39:0] n491;
wire     [47:0] n492;
wire     [55:0] n493;
wire     [63:0] n494;
wire     [71:0] n495;
wire      [7:0] n496;
wire      [7:0] n497;
wire      [7:0] n498;
wire      [7:0] n499;
wire      [7:0] n500;
wire      [7:0] n501;
wire      [7:0] n502;
wire      [7:0] n503;
wire      [7:0] n504;
wire     [15:0] n505;
wire     [23:0] n506;
wire     [31:0] n507;
wire     [39:0] n508;
wire     [47:0] n509;
wire     [55:0] n510;
wire     [63:0] n511;
wire     [71:0] n512;
wire      [7:0] n513;
wire      [7:0] n514;
wire      [7:0] n515;
wire      [7:0] n516;
wire      [7:0] n517;
wire      [7:0] n518;
wire      [7:0] n519;
wire      [7:0] n520;
wire      [7:0] n521;
wire     [15:0] n522;
wire     [23:0] n523;
wire     [31:0] n524;
wire     [39:0] n525;
wire     [47:0] n526;
wire     [55:0] n527;
wire     [63:0] n528;
wire     [71:0] n529;
wire      [7:0] n530;
wire      [7:0] n531;
wire      [7:0] n532;
wire      [7:0] n533;
wire      [7:0] n534;
wire      [7:0] n535;
wire      [7:0] n536;
wire      [7:0] n537;
wire      [7:0] n538;
wire     [15:0] n539;
wire     [23:0] n540;
wire     [31:0] n541;
wire     [39:0] n542;
wire     [47:0] n543;
wire     [55:0] n544;
wire     [63:0] n545;
wire     [71:0] n546;
wire    [143:0] n547;
wire    [215:0] n548;
wire    [287:0] n549;
wire    [359:0] n550;
wire    [431:0] n551;
wire    [503:0] n552;
wire    [575:0] n553;
wire    [647:0] n554;
wire    [647:0] n555;
wire    [647:0] n556;
wire    [647:0] n557;
wire    [647:0] n558;
wire    [647:0] n559;
wire    [647:0] n560;
wire    [647:0] n561;
wire    [647:0] n562;
wire    [647:0] n563;
wire    [647:0] n564;
wire    [647:0] n565;
wire            n566;
wire            n567;
wire            n568;
wire            n569;
wire            n570;
wire            n571;
wire            n572;
wire            n573;
wire            n574;
wire            n575;
wire            n576;
wire            n577;
wire            n578;
wire            n579;
wire            n580;
wire            n581;
wire      [8:0] LB2D_proc_0_addr0;
wire      [7:0] LB2D_proc_0_data0;
wire            n582;
wire            n583;
wire            n584;
wire            n585;
wire            n586;
wire            n587;
wire            n588;
wire            n589;
wire            n590;
wire            n591;
wire            n592;
wire            n593;
wire            n594;
wire            n595;
wire            n596;
wire            n597;
wire      [8:0] LB2D_proc_1_addr0;
wire      [7:0] LB2D_proc_1_data0;
wire            n598;
wire            n599;
wire            n600;
wire      [8:0] LB2D_proc_2_addr0;
wire      [7:0] LB2D_proc_2_data0;
wire            n601;
wire            n602;
wire            n603;
wire      [8:0] LB2D_proc_3_addr0;
wire      [7:0] LB2D_proc_3_data0;
wire            n604;
wire            n605;
wire            n606;
wire      [8:0] LB2D_proc_4_addr0;
wire      [7:0] LB2D_proc_4_data0;
wire            n607;
wire            n608;
wire            n609;
wire      [8:0] LB2D_proc_5_addr0;
wire      [7:0] LB2D_proc_5_data0;
wire            n610;
wire            n611;
wire            n612;
wire      [8:0] LB2D_proc_6_addr0;
wire      [7:0] LB2D_proc_6_data0;
wire            n613;
wire            n614;
wire            n615;
wire      [8:0] LB2D_proc_7_addr0;
wire      [7:0] LB2D_proc_7_data0;
wire            n616;
wire            n617;
wire            n618;
reg      [7:0] LB2D_proc_0[511:0];
reg      [7:0] LB2D_proc_1[511:0];
reg      [7:0] LB2D_proc_2[511:0];
reg      [7:0] LB2D_proc_3[511:0];
reg      [7:0] LB2D_proc_4[511:0];
reg      [7:0] LB2D_proc_5[511:0];
reg      [7:0] LB2D_proc_6[511:0];
reg      [7:0] LB2D_proc_7[511:0];
wire clk;
wire rst;
wire step;
assign n0 =  ( arg_0_TREADY ) == ( 1'd1 )  ;
assign n1 =  ( arg_0_TVALID ) == ( 1'd1 )  ;
assign n2 =  ( n0 ) & ( n1 )  ;
assign n3 =  ( arg_1_TVALID ) == ( 1'd0 )  ;
assign n4 =  ( n2 ) & ( n3 )  ;
assign n5 =  ( arg_0_TVALID ) == ( 1'd0 )  ;
assign n6 =  ( gb_exit_it_1 ) == ( 1'd0 )  ;
assign n7 =  ( stencil_stream_empty ) == ( 1'd0 )  ;
assign n8 =  ( n6 ) & ( n7 )  ;
assign n9 =  ( gb_exit_it_1 ) == ( 1'd1 )  ;
assign n10 =  ( gb_exit_it_8 ) == ( 1'd0 )  ;
assign n11 =  ( n9 ) & ( n10 )  ;
assign n12 =  ( n8 ) | ( n11 )  ;
assign n13 =  ( n5 ) & ( n12 )  ;
assign n14 =  ( slice_stream_empty ) == ( 1'd0 )  ;
assign n15 =  ( LB2D_shift_x ) != ( 9'd488 )  ;
assign n16 =  ( n14 ) & ( n15 )  ;
assign n17 =  ( stencil_stream_full ) == ( 1'd0 )  ;
assign n18 =  ( LB2D_shift_x ) < ( 9'd8 )  ;
assign n19 =  ( n17 ) | ( n18 )  ;
assign n20 =  ( n16 ) & ( n19 )  ;
assign n21 =  ( in_stream_empty ) == ( 1'd0 )  ;
assign n22 =  ( slice_stream_full ) == ( 1'd0 )  ;
assign n23 =  ( LB2D_proc_y ) < ( 10'd8 )  ;
assign n24 =  ( n22 ) | ( n23 )  ;
assign n25 =  ( n21 ) & ( n24 )  ;
assign n26 =  ( arg_1_TREADY ) == ( 1'd0 )  ;
assign n27 =  ( in_stream_full ) == ( 1'd0 )  ;
assign n28 =  ( n26 ) & ( n27 )  ;
assign n29 =  ( LB1D_it_1 ) == ( 1'd0 )  ;
assign n30 =  ( n28 ) & ( n29 )  ;
assign n31 =  ( LB1D_it_1 ) == ( 1'd1 )  ;
assign n32 =  ( n28 ) & ( n31 )  ;
assign n33 =  ( n32 ) ? ( LB1D_uIn ) : ( LB1D_buff ) ;
assign n34 =  ( n30 ) ? ( LB1D_uIn ) : ( n33 ) ;
assign n35 =  ( n25 ) ? ( LB1D_buff ) : ( n34 ) ;
assign n36 =  ( n20 ) ? ( LB1D_buff ) : ( n35 ) ;
assign n37 =  ( n13 ) ? ( LB1D_buff ) : ( n36 ) ;
assign n38 =  ( n4 ) ? ( LB1D_buff ) : ( n37 ) ;
assign n39 =  ( n32 ) ? ( LB1D_in ) : ( LB1D_in ) ;
assign n40 =  ( n30 ) ? ( LB1D_in ) : ( n39 ) ;
assign n41 =  ( n25 ) ? ( LB1D_in ) : ( n40 ) ;
assign n42 =  ( n20 ) ? ( LB1D_in ) : ( n41 ) ;
assign n43 =  ( n13 ) ? ( LB1D_in ) : ( n42 ) ;
assign n44 =  ( n4 ) ? ( LB1D_in ) : ( n43 ) ;
assign n45 =  ( n30 ) ? ( 1'd1 ) : ( LB1D_it_1 ) ;
assign n46 =  ( LB1D_p_cnt ) + ( 19'd1 )  ;
assign n47 =  ( 19'd316224 ) - ( 19'd1 )  ;
assign n48 =  ( LB1D_p_cnt ) == ( n47 )  ;
assign n49 =  ( n48 ) ? ( 19'd0 ) : ( n46 ) ;
assign n50 =  ( n32 ) ? ( n49 ) : ( LB1D_p_cnt ) ;
assign n51 =  ( n30 ) ? ( n46 ) : ( n50 ) ;
assign n52 =  ( n25 ) ? ( LB1D_p_cnt ) : ( n51 ) ;
assign n53 =  ( n20 ) ? ( LB1D_p_cnt ) : ( n52 ) ;
assign n54 =  ( n13 ) ? ( LB1D_p_cnt ) : ( n53 ) ;
assign n55 =  ( n4 ) ? ( LB1D_p_cnt ) : ( n54 ) ;
assign n56 =  ( n32 ) ? ( LB1D_in ) : ( LB1D_uIn ) ;
assign n57 =  ( n30 ) ? ( LB1D_in ) : ( n56 ) ;
assign n58 =  ( n25 ) ? ( LB1D_uIn ) : ( n57 ) ;
assign n59 =  ( n20 ) ? ( LB1D_uIn ) : ( n58 ) ;
assign n60 =  ( n13 ) ? ( LB1D_uIn ) : ( n59 ) ;
assign n61 =  ( LB2D_proc_x ) == ( 9'd488 )  ;
assign n62 =  ( LB2D_proc_w ) == ( 64'd7 )  ;
assign n63 =  ( LB2D_proc_w ) + ( 64'd1 )  ;
assign n64 =  ( n62 ) ? ( 64'd0 ) : ( n63 ) ;
assign n65 =  ( n61 ) ? ( n64 ) : ( LB2D_proc_w ) ;
assign n66 =  ( n32 ) ? ( LB2D_proc_w ) : ( LB2D_proc_w ) ;
assign n67 =  ( n25 ) ? ( n65 ) : ( n66 ) ;
assign n68 =  ( n20 ) ? ( LB2D_proc_w ) : ( n67 ) ;
assign n69 =  ( n13 ) ? ( LB2D_proc_w ) : ( n68 ) ;
assign n70 =  ( n4 ) ? ( LB2D_proc_w ) : ( n69 ) ;
assign n71 =  ( LB2D_proc_x ) + ( 9'd1 )  ;
assign n72 =  ( n61 ) ? ( 9'd1 ) : ( n71 ) ;
assign n73 =  ( n32 ) ? ( LB2D_proc_x ) : ( LB2D_proc_x ) ;
assign n74 =  ( n25 ) ? ( n72 ) : ( n73 ) ;
assign n75 =  ( n20 ) ? ( LB2D_proc_x ) : ( n74 ) ;
assign n76 =  ( n13 ) ? ( LB2D_proc_x ) : ( n75 ) ;
assign n77 =  ( n4 ) ? ( LB2D_proc_x ) : ( n76 ) ;
assign n78 =  ( LB2D_proc_y ) == ( 10'd648 )  ;
assign n79 =  ( LB2D_proc_y ) + ( 10'd1 )  ;
assign n80 =  ( n78 ) ? ( 10'd0 ) : ( n79 ) ;
assign n81 =  ( n61 ) ? ( n80 ) : ( LB2D_proc_y ) ;
assign n82 =  ( n32 ) ? ( LB2D_proc_y ) : ( LB2D_proc_y ) ;
assign n83 =  ( n25 ) ? ( n81 ) : ( n82 ) ;
assign n84 =  ( n20 ) ? ( LB2D_proc_y ) : ( n83 ) ;
assign n85 =  ( n13 ) ? ( LB2D_proc_y ) : ( n84 ) ;
assign n86 =  ( n4 ) ? ( LB2D_proc_y ) : ( n85 ) ;
assign n87 =  ( n32 ) ? ( LB2D_shift_0 ) : ( LB2D_shift_0 ) ;
assign n88 =  ( n25 ) ? ( LB2D_shift_0 ) : ( n87 ) ;
assign n89 =  ( n20 ) ? ( LB2D_shift_1 ) : ( n88 ) ;
assign n90 =  ( n13 ) ? ( LB2D_shift_0 ) : ( n89 ) ;
assign n91 =  ( n4 ) ? ( LB2D_shift_0 ) : ( n90 ) ;
assign n92 =  ( n32 ) ? ( LB2D_shift_1 ) : ( LB2D_shift_1 ) ;
assign n93 =  ( n25 ) ? ( LB2D_shift_1 ) : ( n92 ) ;
assign n94 =  ( n20 ) ? ( LB2D_shift_2 ) : ( n93 ) ;
assign n95 =  ( n13 ) ? ( LB2D_shift_1 ) : ( n94 ) ;
assign n96 =  ( n4 ) ? ( LB2D_shift_1 ) : ( n95 ) ;
assign n97 =  ( n32 ) ? ( LB2D_shift_2 ) : ( LB2D_shift_2 ) ;
assign n98 =  ( n25 ) ? ( LB2D_shift_2 ) : ( n97 ) ;
assign n99 =  ( n20 ) ? ( LB2D_shift_3 ) : ( n98 ) ;
assign n100 =  ( n13 ) ? ( LB2D_shift_2 ) : ( n99 ) ;
assign n101 =  ( n4 ) ? ( LB2D_shift_2 ) : ( n100 ) ;
assign n102 =  ( n32 ) ? ( LB2D_shift_3 ) : ( LB2D_shift_3 ) ;
assign n103 =  ( n25 ) ? ( LB2D_shift_3 ) : ( n102 ) ;
assign n104 =  ( n20 ) ? ( LB2D_shift_4 ) : ( n103 ) ;
assign n105 =  ( n13 ) ? ( LB2D_shift_3 ) : ( n104 ) ;
assign n106 =  ( n4 ) ? ( LB2D_shift_3 ) : ( n105 ) ;
assign n107 =  ( n32 ) ? ( LB2D_shift_4 ) : ( LB2D_shift_4 ) ;
assign n108 =  ( n25 ) ? ( LB2D_shift_4 ) : ( n107 ) ;
assign n109 =  ( n20 ) ? ( LB2D_shift_5 ) : ( n108 ) ;
assign n110 =  ( n13 ) ? ( LB2D_shift_4 ) : ( n109 ) ;
assign n111 =  ( n4 ) ? ( LB2D_shift_4 ) : ( n110 ) ;
assign n112 =  ( n32 ) ? ( LB2D_shift_5 ) : ( LB2D_shift_5 ) ;
assign n113 =  ( n25 ) ? ( LB2D_shift_5 ) : ( n112 ) ;
assign n114 =  ( n20 ) ? ( LB2D_shift_6 ) : ( n113 ) ;
assign n115 =  ( n13 ) ? ( LB2D_shift_5 ) : ( n114 ) ;
assign n116 =  ( n4 ) ? ( LB2D_shift_5 ) : ( n115 ) ;
assign n117 =  ( n32 ) ? ( LB2D_shift_6 ) : ( LB2D_shift_6 ) ;
assign n118 =  ( n25 ) ? ( LB2D_shift_6 ) : ( n117 ) ;
assign n119 =  ( n20 ) ? ( LB2D_shift_7 ) : ( n118 ) ;
assign n120 =  ( n13 ) ? ( LB2D_shift_6 ) : ( n119 ) ;
assign n121 =  ( n4 ) ? ( LB2D_shift_6 ) : ( n120 ) ;
assign n122 =  ( slice_stream_full ) == ( 1'd1 )  ;
assign n123 =  ( n122 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n124 =  ( n32 ) ? ( LB2D_shift_7 ) : ( LB2D_shift_7 ) ;
assign n125 =  ( n25 ) ? ( LB2D_shift_7 ) : ( n124 ) ;
assign n126 =  ( n20 ) ? ( n123 ) : ( n125 ) ;
assign n127 =  ( n13 ) ? ( LB2D_shift_7 ) : ( n126 ) ;
assign n128 =  ( n4 ) ? ( LB2D_shift_7 ) : ( n127 ) ;
assign n129 =  ( LB2D_shift_x ) + ( 9'd1 )  ;
assign n130 =  ( n32 ) ? ( LB2D_shift_x ) : ( LB2D_shift_x ) ;
assign n131 =  ( n25 ) ? ( LB2D_shift_x ) : ( n130 ) ;
assign n132 =  ( n20 ) ? ( n129 ) : ( n131 ) ;
assign n133 =  ( n13 ) ? ( LB2D_shift_x ) : ( n132 ) ;
assign n134 =  ( n4 ) ? ( LB2D_shift_x ) : ( n133 ) ;
assign n135 =  ( LB2D_shift_y ) < ( 10'd640 )  ;
assign n136 =  ( LB2D_shift_x ) < ( 9'd488 )  ;
assign n137 =  ( LB2D_shift_y ) + ( 10'd1 )  ;
assign n138 =  ( n136 ) ? ( LB2D_shift_y ) : ( n137 ) ;
assign n139 =  ( n135 ) ? ( n138 ) : ( 10'd640 ) ;
assign n140 =  ( n32 ) ? ( LB2D_shift_y ) : ( LB2D_shift_y ) ;
assign n141 =  ( n25 ) ? ( LB2D_shift_y ) : ( n140 ) ;
assign n142 =  ( n20 ) ? ( n139 ) : ( n141 ) ;
assign n143 =  ( n13 ) ? ( LB2D_shift_y ) : ( n142 ) ;
assign n144 =  ( n4 ) ? ( LB2D_shift_y ) : ( n143 ) ;
assign n145 =  ( stencil_stream_full ) == ( 1'd1 )  ;
assign n146 =  ( n145 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_0 ) ;
assign n147 = gb_fun(n146) ;
assign n148 =  ( n32 ) ? ( arg_0_TDATA ) : ( arg_0_TDATA ) ;
assign n149 =  ( n25 ) ? ( arg_0_TDATA ) : ( n148 ) ;
assign n150 =  ( n20 ) ? ( arg_0_TDATA ) : ( n149 ) ;
assign n151 =  ( n13 ) ? ( n147 ) : ( n150 ) ;
assign n152 =  ( n4 ) ? ( arg_0_TDATA ) : ( n151 ) ;
assign n153 =  ( gb_pp_it_8 ) == ( 1'd1 )  ;
assign n154 =  ( n153 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n155 =  ( n32 ) ? ( arg_0_TVALID ) : ( arg_0_TVALID ) ;
assign n156 =  ( n25 ) ? ( arg_0_TVALID ) : ( n155 ) ;
assign n157 =  ( n20 ) ? ( arg_0_TVALID ) : ( n156 ) ;
assign n158 =  ( n13 ) ? ( n154 ) : ( n157 ) ;
assign n159 =  ( n4 ) ? ( 1'd0 ) : ( n158 ) ;
assign n160 =  ( n32 ) ? ( 1'd1 ) : ( arg_1_TREADY ) ;
assign n161 =  ( n30 ) ? ( 1'd1 ) : ( n160 ) ;
assign n162 =  ( n25 ) ? ( arg_1_TREADY ) : ( n161 ) ;
assign n163 =  ( n20 ) ? ( arg_1_TREADY ) : ( n162 ) ;
assign n164 =  ( n13 ) ? ( arg_1_TREADY ) : ( n163 ) ;
assign n165 =  ( n4 ) ? ( arg_1_TREADY ) : ( n164 ) ;
assign n166 =  ( gb_p_cnt ) + ( 19'd1 )  ;
assign n167 =  ( n166 ) == ( 19'd307200 )  ;
assign n168 =  ( n167 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n169 =  ( n32 ) ? ( gb_exit_it_1 ) : ( gb_exit_it_1 ) ;
assign n170 =  ( n25 ) ? ( gb_exit_it_1 ) : ( n169 ) ;
assign n171 =  ( n20 ) ? ( gb_exit_it_1 ) : ( n170 ) ;
assign n172 =  ( n13 ) ? ( n168 ) : ( n171 ) ;
assign n173 =  ( n4 ) ? ( gb_exit_it_1 ) : ( n172 ) ;
assign n174 =  ( n32 ) ? ( gb_exit_it_2 ) : ( gb_exit_it_2 ) ;
assign n175 =  ( n25 ) ? ( gb_exit_it_2 ) : ( n174 ) ;
assign n176 =  ( n20 ) ? ( gb_exit_it_2 ) : ( n175 ) ;
assign n177 =  ( n13 ) ? ( gb_exit_it_1 ) : ( n176 ) ;
assign n178 =  ( n4 ) ? ( gb_exit_it_2 ) : ( n177 ) ;
assign n179 =  ( n32 ) ? ( gb_exit_it_3 ) : ( gb_exit_it_3 ) ;
assign n180 =  ( n25 ) ? ( gb_exit_it_3 ) : ( n179 ) ;
assign n181 =  ( n20 ) ? ( gb_exit_it_3 ) : ( n180 ) ;
assign n182 =  ( n13 ) ? ( gb_exit_it_2 ) : ( n181 ) ;
assign n183 =  ( n4 ) ? ( gb_exit_it_3 ) : ( n182 ) ;
assign n184 =  ( n32 ) ? ( gb_exit_it_4 ) : ( gb_exit_it_4 ) ;
assign n185 =  ( n25 ) ? ( gb_exit_it_4 ) : ( n184 ) ;
assign n186 =  ( n20 ) ? ( gb_exit_it_4 ) : ( n185 ) ;
assign n187 =  ( n13 ) ? ( gb_exit_it_3 ) : ( n186 ) ;
assign n188 =  ( n4 ) ? ( gb_exit_it_4 ) : ( n187 ) ;
assign n189 =  ( n32 ) ? ( gb_exit_it_5 ) : ( gb_exit_it_5 ) ;
assign n190 =  ( n25 ) ? ( gb_exit_it_5 ) : ( n189 ) ;
assign n191 =  ( n20 ) ? ( gb_exit_it_5 ) : ( n190 ) ;
assign n192 =  ( n13 ) ? ( gb_exit_it_4 ) : ( n191 ) ;
assign n193 =  ( n4 ) ? ( gb_exit_it_5 ) : ( n192 ) ;
assign n194 =  ( n32 ) ? ( gb_exit_it_6 ) : ( gb_exit_it_6 ) ;
assign n195 =  ( n25 ) ? ( gb_exit_it_6 ) : ( n194 ) ;
assign n196 =  ( n20 ) ? ( gb_exit_it_6 ) : ( n195 ) ;
assign n197 =  ( n13 ) ? ( gb_exit_it_5 ) : ( n196 ) ;
assign n198 =  ( n4 ) ? ( gb_exit_it_6 ) : ( n197 ) ;
assign n199 =  ( n32 ) ? ( gb_exit_it_7 ) : ( gb_exit_it_7 ) ;
assign n200 =  ( n25 ) ? ( gb_exit_it_7 ) : ( n199 ) ;
assign n201 =  ( n20 ) ? ( gb_exit_it_7 ) : ( n200 ) ;
assign n202 =  ( n13 ) ? ( gb_exit_it_6 ) : ( n201 ) ;
assign n203 =  ( n4 ) ? ( gb_exit_it_7 ) : ( n202 ) ;
assign n204 =  ( n32 ) ? ( gb_exit_it_8 ) : ( gb_exit_it_8 ) ;
assign n205 =  ( n25 ) ? ( gb_exit_it_8 ) : ( n204 ) ;
assign n206 =  ( n20 ) ? ( gb_exit_it_8 ) : ( n205 ) ;
assign n207 =  ( n13 ) ? ( gb_exit_it_7 ) : ( n206 ) ;
assign n208 =  ( n4 ) ? ( gb_exit_it_8 ) : ( n207 ) ;
assign n209 =  ( gb_p_cnt ) < ( 19'd307200 )  ;
assign n210 =  ( n209 ) ? ( n166 ) : ( 19'd307200 ) ;
assign n211 =  ( n32 ) ? ( gb_p_cnt ) : ( gb_p_cnt ) ;
assign n212 =  ( n25 ) ? ( gb_p_cnt ) : ( n211 ) ;
assign n213 =  ( n20 ) ? ( gb_p_cnt ) : ( n212 ) ;
assign n214 =  ( n13 ) ? ( n210 ) : ( n213 ) ;
assign n215 =  ( n4 ) ? ( gb_p_cnt ) : ( n214 ) ;
assign n216 =  ( n32 ) ? ( gb_pp_it_1 ) : ( gb_pp_it_1 ) ;
assign n217 =  ( n25 ) ? ( gb_pp_it_1 ) : ( n216 ) ;
assign n218 =  ( n20 ) ? ( gb_pp_it_1 ) : ( n217 ) ;
assign n219 =  ( n13 ) ? ( 1'd1 ) : ( n218 ) ;
assign n220 =  ( n4 ) ? ( gb_pp_it_1 ) : ( n219 ) ;
assign n221 =  ( n32 ) ? ( gb_pp_it_2 ) : ( gb_pp_it_2 ) ;
assign n222 =  ( n25 ) ? ( gb_pp_it_2 ) : ( n221 ) ;
assign n223 =  ( n20 ) ? ( gb_pp_it_2 ) : ( n222 ) ;
assign n224 =  ( n13 ) ? ( gb_pp_it_1 ) : ( n223 ) ;
assign n225 =  ( n4 ) ? ( gb_pp_it_2 ) : ( n224 ) ;
assign n226 =  ( n32 ) ? ( gb_pp_it_3 ) : ( gb_pp_it_3 ) ;
assign n227 =  ( n25 ) ? ( gb_pp_it_3 ) : ( n226 ) ;
assign n228 =  ( n20 ) ? ( gb_pp_it_3 ) : ( n227 ) ;
assign n229 =  ( n13 ) ? ( gb_pp_it_2 ) : ( n228 ) ;
assign n230 =  ( n4 ) ? ( gb_pp_it_3 ) : ( n229 ) ;
assign n231 =  ( n32 ) ? ( gb_pp_it_4 ) : ( gb_pp_it_4 ) ;
assign n232 =  ( n25 ) ? ( gb_pp_it_4 ) : ( n231 ) ;
assign n233 =  ( n20 ) ? ( gb_pp_it_4 ) : ( n232 ) ;
assign n234 =  ( n13 ) ? ( gb_pp_it_3 ) : ( n233 ) ;
assign n235 =  ( n4 ) ? ( gb_pp_it_4 ) : ( n234 ) ;
assign n236 =  ( n32 ) ? ( gb_pp_it_5 ) : ( gb_pp_it_5 ) ;
assign n237 =  ( n25 ) ? ( gb_pp_it_5 ) : ( n236 ) ;
assign n238 =  ( n20 ) ? ( gb_pp_it_5 ) : ( n237 ) ;
assign n239 =  ( n13 ) ? ( gb_pp_it_4 ) : ( n238 ) ;
assign n240 =  ( n4 ) ? ( gb_pp_it_5 ) : ( n239 ) ;
assign n241 =  ( n32 ) ? ( gb_pp_it_6 ) : ( gb_pp_it_6 ) ;
assign n242 =  ( n25 ) ? ( gb_pp_it_6 ) : ( n241 ) ;
assign n243 =  ( n20 ) ? ( gb_pp_it_6 ) : ( n242 ) ;
assign n244 =  ( n13 ) ? ( gb_pp_it_5 ) : ( n243 ) ;
assign n245 =  ( n4 ) ? ( gb_pp_it_6 ) : ( n244 ) ;
assign n246 =  ( n32 ) ? ( gb_pp_it_7 ) : ( gb_pp_it_7 ) ;
assign n247 =  ( n25 ) ? ( gb_pp_it_7 ) : ( n246 ) ;
assign n248 =  ( n20 ) ? ( gb_pp_it_7 ) : ( n247 ) ;
assign n249 =  ( n13 ) ? ( gb_pp_it_6 ) : ( n248 ) ;
assign n250 =  ( n4 ) ? ( gb_pp_it_7 ) : ( n249 ) ;
assign n251 =  ( n32 ) ? ( gb_pp_it_8 ) : ( gb_pp_it_8 ) ;
assign n252 =  ( n25 ) ? ( gb_pp_it_8 ) : ( n251 ) ;
assign n253 =  ( n20 ) ? ( gb_pp_it_8 ) : ( n252 ) ;
assign n254 =  ( n13 ) ? ( gb_pp_it_7 ) : ( n253 ) ;
assign n255 =  ( n4 ) ? ( gb_pp_it_8 ) : ( n254 ) ;
assign n256 =  ( n32 ) ? ( gb_pp_it_9 ) : ( gb_pp_it_9 ) ;
assign n257 =  ( n25 ) ? ( gb_pp_it_9 ) : ( n256 ) ;
assign n258 =  ( n20 ) ? ( gb_pp_it_9 ) : ( n257 ) ;
assign n259 =  ( n13 ) ? ( gb_pp_it_8 ) : ( n258 ) ;
assign n260 =  ( n4 ) ? ( gb_pp_it_9 ) : ( n259 ) ;
assign n261 =  ( n32 ) ? ( LB1D_buff ) : ( in_stream_buff_0 ) ;
assign n262 =  ( n25 ) ? ( in_stream_buff_0 ) : ( n261 ) ;
assign n263 =  ( n20 ) ? ( in_stream_buff_0 ) : ( n262 ) ;
assign n264 =  ( n13 ) ? ( in_stream_buff_0 ) : ( n263 ) ;
assign n265 =  ( n4 ) ? ( in_stream_buff_0 ) : ( n264 ) ;
assign n266 =  ( n32 ) ? ( in_stream_buff_0 ) : ( in_stream_buff_1 ) ;
assign n267 =  ( n25 ) ? ( in_stream_buff_1 ) : ( n266 ) ;
assign n268 =  ( n20 ) ? ( in_stream_buff_1 ) : ( n267 ) ;
assign n269 =  ( n13 ) ? ( in_stream_buff_1 ) : ( n268 ) ;
assign n270 =  ( n4 ) ? ( in_stream_buff_1 ) : ( n269 ) ;
assign n271 =  ( in_stream_full ) == ( 1'd1 )  ;
assign n272 =  ( n271 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n273 =  ( n32 ) ? ( 1'd0 ) : ( in_stream_empty ) ;
assign n274 =  ( n25 ) ? ( n272 ) : ( n273 ) ;
assign n275 =  ( n20 ) ? ( in_stream_empty ) : ( n274 ) ;
assign n276 =  ( n13 ) ? ( in_stream_empty ) : ( n275 ) ;
assign n277 =  ( n4 ) ? ( in_stream_empty ) : ( n276 ) ;
assign n278 =  ( in_stream_empty ) == ( 1'd1 )  ;
assign n279 =  ( n278 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n280 =  ( n32 ) ? ( n279 ) : ( in_stream_full ) ;
assign n281 =  ( n25 ) ? ( 1'd0 ) : ( n280 ) ;
assign n282 =  ( n20 ) ? ( in_stream_full ) : ( n281 ) ;
assign n283 =  ( n13 ) ? ( in_stream_full ) : ( n282 ) ;
assign n284 =  ( n4 ) ? ( in_stream_full ) : ( n283 ) ;
assign n285 =  ( n271 ) ? ( in_stream_buff_1 ) : ( in_stream_buff_0 ) ;
assign n286 =  ( LB2D_proc_w ) == ( 64'd0 )  ;
assign n287 =  ( LB2D_proc_x ) - ( 9'd1 )  ;
assign n288 =  (  LB2D_proc_7 [ n287 ] )  ;
assign n289 =  ( LB2D_proc_w ) == ( 64'd1 )  ;
assign n290 =  (  LB2D_proc_0 [ n287 ] )  ;
assign n291 =  ( LB2D_proc_w ) == ( 64'd2 )  ;
assign n292 =  (  LB2D_proc_1 [ n287 ] )  ;
assign n293 =  ( LB2D_proc_w ) == ( 64'd3 )  ;
assign n294 =  (  LB2D_proc_2 [ n287 ] )  ;
assign n295 =  ( LB2D_proc_w ) == ( 64'd4 )  ;
assign n296 =  (  LB2D_proc_3 [ n287 ] )  ;
assign n297 =  ( LB2D_proc_w ) == ( 64'd5 )  ;
assign n298 =  (  LB2D_proc_4 [ n287 ] )  ;
assign n299 =  ( LB2D_proc_w ) == ( 64'd6 )  ;
assign n300 =  (  LB2D_proc_5 [ n287 ] )  ;
assign n301 =  (  LB2D_proc_6 [ n287 ] )  ;
assign n302 =  ( n299 ) ? ( n300 ) : ( n301 ) ;
assign n303 =  ( n297 ) ? ( n298 ) : ( n302 ) ;
assign n304 =  ( n295 ) ? ( n296 ) : ( n303 ) ;
assign n305 =  ( n293 ) ? ( n294 ) : ( n304 ) ;
assign n306 =  ( n291 ) ? ( n292 ) : ( n305 ) ;
assign n307 =  ( n289 ) ? ( n290 ) : ( n306 ) ;
assign n308 =  ( n286 ) ? ( n288 ) : ( n307 ) ;
assign n309 =  ( n299 ) ? ( n298 ) : ( n300 ) ;
assign n310 =  ( n297 ) ? ( n296 ) : ( n309 ) ;
assign n311 =  ( n295 ) ? ( n294 ) : ( n310 ) ;
assign n312 =  ( n293 ) ? ( n292 ) : ( n311 ) ;
assign n313 =  ( n291 ) ? ( n290 ) : ( n312 ) ;
assign n314 =  ( n289 ) ? ( n288 ) : ( n313 ) ;
assign n315 =  ( n286 ) ? ( n301 ) : ( n314 ) ;
assign n316 =  ( n299 ) ? ( n296 ) : ( n298 ) ;
assign n317 =  ( n297 ) ? ( n294 ) : ( n316 ) ;
assign n318 =  ( n295 ) ? ( n292 ) : ( n317 ) ;
assign n319 =  ( n293 ) ? ( n290 ) : ( n318 ) ;
assign n320 =  ( n291 ) ? ( n288 ) : ( n319 ) ;
assign n321 =  ( n289 ) ? ( n301 ) : ( n320 ) ;
assign n322 =  ( n286 ) ? ( n300 ) : ( n321 ) ;
assign n323 =  ( n299 ) ? ( n294 ) : ( n296 ) ;
assign n324 =  ( n297 ) ? ( n292 ) : ( n323 ) ;
assign n325 =  ( n295 ) ? ( n290 ) : ( n324 ) ;
assign n326 =  ( n293 ) ? ( n288 ) : ( n325 ) ;
assign n327 =  ( n291 ) ? ( n301 ) : ( n326 ) ;
assign n328 =  ( n289 ) ? ( n300 ) : ( n327 ) ;
assign n329 =  ( n286 ) ? ( n298 ) : ( n328 ) ;
assign n330 =  ( n299 ) ? ( n292 ) : ( n294 ) ;
assign n331 =  ( n297 ) ? ( n290 ) : ( n330 ) ;
assign n332 =  ( n295 ) ? ( n288 ) : ( n331 ) ;
assign n333 =  ( n293 ) ? ( n301 ) : ( n332 ) ;
assign n334 =  ( n291 ) ? ( n300 ) : ( n333 ) ;
assign n335 =  ( n289 ) ? ( n298 ) : ( n334 ) ;
assign n336 =  ( n286 ) ? ( n296 ) : ( n335 ) ;
assign n337 =  ( n299 ) ? ( n290 ) : ( n292 ) ;
assign n338 =  ( n297 ) ? ( n288 ) : ( n337 ) ;
assign n339 =  ( n295 ) ? ( n301 ) : ( n338 ) ;
assign n340 =  ( n293 ) ? ( n300 ) : ( n339 ) ;
assign n341 =  ( n291 ) ? ( n298 ) : ( n340 ) ;
assign n342 =  ( n289 ) ? ( n296 ) : ( n341 ) ;
assign n343 =  ( n286 ) ? ( n294 ) : ( n342 ) ;
assign n344 =  ( n299 ) ? ( n288 ) : ( n290 ) ;
assign n345 =  ( n297 ) ? ( n301 ) : ( n344 ) ;
assign n346 =  ( n295 ) ? ( n300 ) : ( n345 ) ;
assign n347 =  ( n293 ) ? ( n298 ) : ( n346 ) ;
assign n348 =  ( n291 ) ? ( n296 ) : ( n347 ) ;
assign n349 =  ( n289 ) ? ( n294 ) : ( n348 ) ;
assign n350 =  ( n286 ) ? ( n292 ) : ( n349 ) ;
assign n351 =  ( n299 ) ? ( n301 ) : ( n288 ) ;
assign n352 =  ( n297 ) ? ( n300 ) : ( n351 ) ;
assign n353 =  ( n295 ) ? ( n298 ) : ( n352 ) ;
assign n354 =  ( n293 ) ? ( n296 ) : ( n353 ) ;
assign n355 =  ( n291 ) ? ( n294 ) : ( n354 ) ;
assign n356 =  ( n289 ) ? ( n292 ) : ( n355 ) ;
assign n357 =  ( n286 ) ? ( n290 ) : ( n356 ) ;
assign n358 =  { ( n350 ) , ( n357 ) }  ;
assign n359 =  { ( n343 ) , ( n358 ) }  ;
assign n360 =  { ( n336 ) , ( n359 ) }  ;
assign n361 =  { ( n329 ) , ( n360 ) }  ;
assign n362 =  { ( n322 ) , ( n361 ) }  ;
assign n363 =  { ( n315 ) , ( n362 ) }  ;
assign n364 =  { ( n308 ) , ( n363 ) }  ;
assign n365 =  { ( n285 ) , ( n364 ) }  ;
assign n366 =  ( n23 ) ? ( slice_stream_buff_0 ) : ( n365 ) ;
assign n367 =  ( n32 ) ? ( slice_stream_buff_0 ) : ( slice_stream_buff_0 ) ;
assign n368 =  ( n25 ) ? ( n366 ) : ( n367 ) ;
assign n369 =  ( n20 ) ? ( slice_stream_buff_0 ) : ( n368 ) ;
assign n370 =  ( n13 ) ? ( slice_stream_buff_0 ) : ( n369 ) ;
assign n371 =  ( n4 ) ? ( slice_stream_buff_0 ) : ( n370 ) ;
assign n372 =  ( n23 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n373 =  ( n32 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_1 ) ;
assign n374 =  ( n25 ) ? ( n372 ) : ( n373 ) ;
assign n375 =  ( n20 ) ? ( slice_stream_buff_1 ) : ( n374 ) ;
assign n376 =  ( n13 ) ? ( slice_stream_buff_1 ) : ( n375 ) ;
assign n377 =  ( n4 ) ? ( slice_stream_buff_1 ) : ( n376 ) ;
assign n378 =  ( n122 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n379 =  ( n23 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n380 =  ( n32 ) ? ( slice_stream_empty ) : ( slice_stream_empty ) ;
assign n381 =  ( n25 ) ? ( n379 ) : ( n380 ) ;
assign n382 =  ( n20 ) ? ( n378 ) : ( n381 ) ;
assign n383 =  ( n13 ) ? ( slice_stream_empty ) : ( n382 ) ;
assign n384 =  ( n4 ) ? ( slice_stream_empty ) : ( n383 ) ;
assign n385 =  ( slice_stream_empty ) == ( 1'd1 )  ;
assign n386 =  ( n385 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n387 =  ( n23 ) ? ( 1'd0 ) : ( n386 ) ;
assign n388 =  ( n32 ) ? ( slice_stream_full ) : ( slice_stream_full ) ;
assign n389 =  ( n25 ) ? ( n387 ) : ( n388 ) ;
assign n390 =  ( n20 ) ? ( 1'd0 ) : ( n389 ) ;
assign n391 =  ( n13 ) ? ( slice_stream_full ) : ( n390 ) ;
assign n392 =  ( n4 ) ? ( slice_stream_full ) : ( n391 ) ;
assign n393 =  ( LB2D_shift_x ) >= ( 9'd8 )  ;
assign n394 = n123[71:64] ;
assign n395 = LB2D_shift_7[71:64] ;
assign n396 = LB2D_shift_6[71:64] ;
assign n397 = LB2D_shift_5[71:64] ;
assign n398 = LB2D_shift_4[71:64] ;
assign n399 = LB2D_shift_3[71:64] ;
assign n400 = LB2D_shift_2[71:64] ;
assign n401 = LB2D_shift_1[71:64] ;
assign n402 = LB2D_shift_0[71:64] ;
assign n403 =  { ( n401 ) , ( n402 ) }  ;
assign n404 =  { ( n400 ) , ( n403 ) }  ;
assign n405 =  { ( n399 ) , ( n404 ) }  ;
assign n406 =  { ( n398 ) , ( n405 ) }  ;
assign n407 =  { ( n397 ) , ( n406 ) }  ;
assign n408 =  { ( n396 ) , ( n407 ) }  ;
assign n409 =  { ( n395 ) , ( n408 ) }  ;
assign n410 =  { ( n394 ) , ( n409 ) }  ;
assign n411 = n123[63:56] ;
assign n412 = LB2D_shift_7[63:56] ;
assign n413 = LB2D_shift_6[63:56] ;
assign n414 = LB2D_shift_5[63:56] ;
assign n415 = LB2D_shift_4[63:56] ;
assign n416 = LB2D_shift_3[63:56] ;
assign n417 = LB2D_shift_2[63:56] ;
assign n418 = LB2D_shift_1[63:56] ;
assign n419 = LB2D_shift_0[63:56] ;
assign n420 =  { ( n418 ) , ( n419 ) }  ;
assign n421 =  { ( n417 ) , ( n420 ) }  ;
assign n422 =  { ( n416 ) , ( n421 ) }  ;
assign n423 =  { ( n415 ) , ( n422 ) }  ;
assign n424 =  { ( n414 ) , ( n423 ) }  ;
assign n425 =  { ( n413 ) , ( n424 ) }  ;
assign n426 =  { ( n412 ) , ( n425 ) }  ;
assign n427 =  { ( n411 ) , ( n426 ) }  ;
assign n428 = n123[55:48] ;
assign n429 = LB2D_shift_7[55:48] ;
assign n430 = LB2D_shift_6[55:48] ;
assign n431 = LB2D_shift_5[55:48] ;
assign n432 = LB2D_shift_4[55:48] ;
assign n433 = LB2D_shift_3[55:48] ;
assign n434 = LB2D_shift_2[55:48] ;
assign n435 = LB2D_shift_1[55:48] ;
assign n436 = LB2D_shift_0[55:48] ;
assign n437 =  { ( n435 ) , ( n436 ) }  ;
assign n438 =  { ( n434 ) , ( n437 ) }  ;
assign n439 =  { ( n433 ) , ( n438 ) }  ;
assign n440 =  { ( n432 ) , ( n439 ) }  ;
assign n441 =  { ( n431 ) , ( n440 ) }  ;
assign n442 =  { ( n430 ) , ( n441 ) }  ;
assign n443 =  { ( n429 ) , ( n442 ) }  ;
assign n444 =  { ( n428 ) , ( n443 ) }  ;
assign n445 = n123[47:40] ;
assign n446 = LB2D_shift_7[47:40] ;
assign n447 = LB2D_shift_6[47:40] ;
assign n448 = LB2D_shift_5[47:40] ;
assign n449 = LB2D_shift_4[47:40] ;
assign n450 = LB2D_shift_3[47:40] ;
assign n451 = LB2D_shift_2[47:40] ;
assign n452 = LB2D_shift_1[47:40] ;
assign n453 = LB2D_shift_0[47:40] ;
assign n454 =  { ( n452 ) , ( n453 ) }  ;
assign n455 =  { ( n451 ) , ( n454 ) }  ;
assign n456 =  { ( n450 ) , ( n455 ) }  ;
assign n457 =  { ( n449 ) , ( n456 ) }  ;
assign n458 =  { ( n448 ) , ( n457 ) }  ;
assign n459 =  { ( n447 ) , ( n458 ) }  ;
assign n460 =  { ( n446 ) , ( n459 ) }  ;
assign n461 =  { ( n445 ) , ( n460 ) }  ;
assign n462 = n123[39:32] ;
assign n463 = LB2D_shift_7[39:32] ;
assign n464 = LB2D_shift_6[39:32] ;
assign n465 = LB2D_shift_5[39:32] ;
assign n466 = LB2D_shift_4[39:32] ;
assign n467 = LB2D_shift_3[39:32] ;
assign n468 = LB2D_shift_2[39:32] ;
assign n469 = LB2D_shift_1[39:32] ;
assign n470 = LB2D_shift_0[39:32] ;
assign n471 =  { ( n469 ) , ( n470 ) }  ;
assign n472 =  { ( n468 ) , ( n471 ) }  ;
assign n473 =  { ( n467 ) , ( n472 ) }  ;
assign n474 =  { ( n466 ) , ( n473 ) }  ;
assign n475 =  { ( n465 ) , ( n474 ) }  ;
assign n476 =  { ( n464 ) , ( n475 ) }  ;
assign n477 =  { ( n463 ) , ( n476 ) }  ;
assign n478 =  { ( n462 ) , ( n477 ) }  ;
assign n479 = n123[31:24] ;
assign n480 = LB2D_shift_7[31:24] ;
assign n481 = LB2D_shift_6[31:24] ;
assign n482 = LB2D_shift_5[31:24] ;
assign n483 = LB2D_shift_4[31:24] ;
assign n484 = LB2D_shift_3[31:24] ;
assign n485 = LB2D_shift_2[31:24] ;
assign n486 = LB2D_shift_1[31:24] ;
assign n487 = LB2D_shift_0[31:24] ;
assign n488 =  { ( n486 ) , ( n487 ) }  ;
assign n489 =  { ( n485 ) , ( n488 ) }  ;
assign n490 =  { ( n484 ) , ( n489 ) }  ;
assign n491 =  { ( n483 ) , ( n490 ) }  ;
assign n492 =  { ( n482 ) , ( n491 ) }  ;
assign n493 =  { ( n481 ) , ( n492 ) }  ;
assign n494 =  { ( n480 ) , ( n493 ) }  ;
assign n495 =  { ( n479 ) , ( n494 ) }  ;
assign n496 = n123[23:16] ;
assign n497 = LB2D_shift_7[23:16] ;
assign n498 = LB2D_shift_6[23:16] ;
assign n499 = LB2D_shift_5[23:16] ;
assign n500 = LB2D_shift_4[23:16] ;
assign n501 = LB2D_shift_3[23:16] ;
assign n502 = LB2D_shift_2[23:16] ;
assign n503 = LB2D_shift_1[23:16] ;
assign n504 = LB2D_shift_0[23:16] ;
assign n505 =  { ( n503 ) , ( n504 ) }  ;
assign n506 =  { ( n502 ) , ( n505 ) }  ;
assign n507 =  { ( n501 ) , ( n506 ) }  ;
assign n508 =  { ( n500 ) , ( n507 ) }  ;
assign n509 =  { ( n499 ) , ( n508 ) }  ;
assign n510 =  { ( n498 ) , ( n509 ) }  ;
assign n511 =  { ( n497 ) , ( n510 ) }  ;
assign n512 =  { ( n496 ) , ( n511 ) }  ;
assign n513 = n123[15:8] ;
assign n514 = LB2D_shift_7[15:8] ;
assign n515 = LB2D_shift_6[15:8] ;
assign n516 = LB2D_shift_5[15:8] ;
assign n517 = LB2D_shift_4[15:8] ;
assign n518 = LB2D_shift_3[15:8] ;
assign n519 = LB2D_shift_2[15:8] ;
assign n520 = LB2D_shift_1[15:8] ;
assign n521 = LB2D_shift_0[15:8] ;
assign n522 =  { ( n520 ) , ( n521 ) }  ;
assign n523 =  { ( n519 ) , ( n522 ) }  ;
assign n524 =  { ( n518 ) , ( n523 ) }  ;
assign n525 =  { ( n517 ) , ( n524 ) }  ;
assign n526 =  { ( n516 ) , ( n525 ) }  ;
assign n527 =  { ( n515 ) , ( n526 ) }  ;
assign n528 =  { ( n514 ) , ( n527 ) }  ;
assign n529 =  { ( n513 ) , ( n528 ) }  ;
assign n530 = n123[7:0] ;
assign n531 = LB2D_shift_7[7:0] ;
assign n532 = LB2D_shift_6[7:0] ;
assign n533 = LB2D_shift_5[7:0] ;
assign n534 = LB2D_shift_4[7:0] ;
assign n535 = LB2D_shift_3[7:0] ;
assign n536 = LB2D_shift_2[7:0] ;
assign n537 = LB2D_shift_1[7:0] ;
assign n538 = LB2D_shift_0[7:0] ;
assign n539 =  { ( n537 ) , ( n538 ) }  ;
assign n540 =  { ( n536 ) , ( n539 ) }  ;
assign n541 =  { ( n535 ) , ( n540 ) }  ;
assign n542 =  { ( n534 ) , ( n541 ) }  ;
assign n543 =  { ( n533 ) , ( n542 ) }  ;
assign n544 =  { ( n532 ) , ( n543 ) }  ;
assign n545 =  { ( n531 ) , ( n544 ) }  ;
assign n546 =  { ( n530 ) , ( n545 ) }  ;
assign n547 =  { ( n529 ) , ( n546 ) }  ;
assign n548 =  { ( n512 ) , ( n547 ) }  ;
assign n549 =  { ( n495 ) , ( n548 ) }  ;
assign n550 =  { ( n478 ) , ( n549 ) }  ;
assign n551 =  { ( n461 ) , ( n550 ) }  ;
assign n552 =  { ( n444 ) , ( n551 ) }  ;
assign n553 =  { ( n427 ) , ( n552 ) }  ;
assign n554 =  { ( n410 ) , ( n553 ) }  ;
assign n555 =  ( n393 ) ? ( n554 ) : ( stencil_stream_buff_0 ) ;
assign n556 =  ( n32 ) ? ( stencil_stream_buff_0 ) : ( stencil_stream_buff_0 ) ;
assign n557 =  ( n25 ) ? ( stencil_stream_buff_0 ) : ( n556 ) ;
assign n558 =  ( n20 ) ? ( n555 ) : ( n557 ) ;
assign n559 =  ( n13 ) ? ( stencil_stream_buff_0 ) : ( n558 ) ;
assign n560 =  ( n4 ) ? ( stencil_stream_buff_0 ) : ( n559 ) ;
assign n561 =  ( n32 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_1 ) ;
assign n562 =  ( n25 ) ? ( stencil_stream_buff_1 ) : ( n561 ) ;
assign n563 =  ( n20 ) ? ( stencil_stream_buff_0 ) : ( n562 ) ;
assign n564 =  ( n13 ) ? ( stencil_stream_buff_1 ) : ( n563 ) ;
assign n565 =  ( n4 ) ? ( stencil_stream_buff_1 ) : ( n564 ) ;
assign n566 =  ( n145 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n567 =  ( n18 ) ? ( stencil_stream_empty ) : ( 1'd0 ) ;
assign n568 =  ( n32 ) ? ( stencil_stream_empty ) : ( stencil_stream_empty ) ;
assign n569 =  ( n25 ) ? ( stencil_stream_empty ) : ( n568 ) ;
assign n570 =  ( n20 ) ? ( n567 ) : ( n569 ) ;
assign n571 =  ( n13 ) ? ( n566 ) : ( n570 ) ;
assign n572 =  ( n4 ) ? ( stencil_stream_empty ) : ( n571 ) ;
assign n573 =  ( n9 ) ? ( 1'd0 ) : ( 1'd0 ) ;
assign n574 =  ( stencil_stream_empty ) == ( 1'd1 )  ;
assign n575 =  ( n574 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n576 =  ( n18 ) ? ( stencil_stream_full ) : ( n575 ) ;
assign n577 =  ( n32 ) ? ( stencil_stream_full ) : ( stencil_stream_full ) ;
assign n578 =  ( n25 ) ? ( stencil_stream_full ) : ( n577 ) ;
assign n579 =  ( n20 ) ? ( n576 ) : ( n578 ) ;
assign n580 =  ( n13 ) ? ( n573 ) : ( n579 ) ;
assign n581 =  ( n4 ) ? ( stencil_stream_full ) : ( n580 ) ;
assign n582 = ~ ( n4 ) ;
assign n583 = ~ ( n13 ) ;
assign n584 =  ( n582 ) & ( n583 )  ;
assign n585 = ~ ( n20 ) ;
assign n586 =  ( n584 ) & ( n585 )  ;
assign n587 = ~ ( n25 ) ;
assign n588 =  ( n586 ) & ( n587 )  ;
assign n589 = ~ ( n32 ) ;
assign n590 =  ( n588 ) & ( n589 )  ;
assign n591 =  ( n588 ) & ( n32 )  ;
assign n592 =  ( n586 ) & ( n25 )  ;
assign n593 = ~ ( n286 ) ;
assign n594 =  ( n592 ) & ( n593 )  ;
assign n595 =  ( n592 ) & ( n286 )  ;
assign n596 =  ( n584 ) & ( n20 )  ;
assign n597 =  ( n582 ) & ( n13 )  ;
assign LB2D_proc_0_addr0 = n595 ? (n287) : (0);
assign LB2D_proc_0_data0 = n595 ? (n285) : (LB2D_proc_0[0]);
assign n598 = ~ ( n289 ) ;
assign n599 =  ( n592 ) & ( n598 )  ;
assign n600 =  ( n592 ) & ( n289 )  ;
assign LB2D_proc_1_addr0 = n600 ? (n287) : (0);
assign LB2D_proc_1_data0 = n600 ? (n285) : (LB2D_proc_1[0]);
assign n601 = ~ ( n291 ) ;
assign n602 =  ( n592 ) & ( n601 )  ;
assign n603 =  ( n592 ) & ( n291 )  ;
assign LB2D_proc_2_addr0 = n603 ? (n287) : (0);
assign LB2D_proc_2_data0 = n603 ? (n285) : (LB2D_proc_2[0]);
assign n604 = ~ ( n293 ) ;
assign n605 =  ( n592 ) & ( n604 )  ;
assign n606 =  ( n592 ) & ( n293 )  ;
assign LB2D_proc_3_addr0 = n606 ? (n287) : (0);
assign LB2D_proc_3_data0 = n606 ? (n285) : (LB2D_proc_3[0]);
assign n607 = ~ ( n295 ) ;
assign n608 =  ( n592 ) & ( n607 )  ;
assign n609 =  ( n592 ) & ( n295 )  ;
assign LB2D_proc_4_addr0 = n609 ? (n287) : (0);
assign LB2D_proc_4_data0 = n609 ? (n285) : (LB2D_proc_4[0]);
assign n610 = ~ ( n297 ) ;
assign n611 =  ( n592 ) & ( n610 )  ;
assign n612 =  ( n592 ) & ( n297 )  ;
assign LB2D_proc_5_addr0 = n612 ? (n287) : (0);
assign LB2D_proc_5_data0 = n612 ? (n285) : (LB2D_proc_5[0]);
assign n613 = ~ ( n299 ) ;
assign n614 =  ( n592 ) & ( n613 )  ;
assign n615 =  ( n592 ) & ( n299 )  ;
assign LB2D_proc_6_addr0 = n615 ? (n287) : (0);
assign LB2D_proc_6_data0 = n615 ? (n285) : (LB2D_proc_6[0]);
assign n616 = ~ ( n62 ) ;
assign n617 =  ( n592 ) & ( n616 )  ;
assign n618 =  ( n592 ) & ( n62 )  ;
assign LB2D_proc_7_addr0 = n618 ? (n287) : (0);
assign LB2D_proc_7_data0 = n618 ? (n285) : (LB2D_proc_7[0]);
/*
function [7:0] gb_fun ;
input [647:0] arg0;
    begin
//TODO: Add the specific function HERE.    end
endfunction
*/

always @(posedge clk) begin
   if(rst) begin
       LB1D_buff <= LB1D_buff;
       LB1D_in <= LB1D_in;
       LB1D_it_1 <= LB1D_it_1;
       LB1D_p_cnt <= LB1D_p_cnt;
       LB1D_uIn <= LB1D_uIn;
       LB2D_proc_w <= LB2D_proc_w;
       LB2D_proc_x <= LB2D_proc_x;
       LB2D_proc_y <= LB2D_proc_y;
       LB2D_shift_0 <= LB2D_shift_0;
       LB2D_shift_1 <= LB2D_shift_1;
       LB2D_shift_2 <= LB2D_shift_2;
       LB2D_shift_3 <= LB2D_shift_3;
       LB2D_shift_4 <= LB2D_shift_4;
       LB2D_shift_5 <= LB2D_shift_5;
       LB2D_shift_6 <= LB2D_shift_6;
       LB2D_shift_7 <= LB2D_shift_7;
       LB2D_shift_x <= LB2D_shift_x;
       LB2D_shift_y <= LB2D_shift_y;
       arg_0_TDATA <= arg_0_TDATA;
       arg_0_TVALID <= arg_0_TVALID;
       arg_1_TREADY <= arg_1_TREADY;
       gb_exit_it_1 <= gb_exit_it_1;
       gb_exit_it_2 <= gb_exit_it_2;
       gb_exit_it_3 <= gb_exit_it_3;
       gb_exit_it_4 <= gb_exit_it_4;
       gb_exit_it_5 <= gb_exit_it_5;
       gb_exit_it_6 <= gb_exit_it_6;
       gb_exit_it_7 <= gb_exit_it_7;
       gb_exit_it_8 <= gb_exit_it_8;
       gb_p_cnt <= gb_p_cnt;
       gb_pp_it_1 <= gb_pp_it_1;
       gb_pp_it_2 <= gb_pp_it_2;
       gb_pp_it_3 <= gb_pp_it_3;
       gb_pp_it_4 <= gb_pp_it_4;
       gb_pp_it_5 <= gb_pp_it_5;
       gb_pp_it_6 <= gb_pp_it_6;
       gb_pp_it_7 <= gb_pp_it_7;
       gb_pp_it_8 <= gb_pp_it_8;
       gb_pp_it_9 <= gb_pp_it_9;
       in_stream_buff_0 <= in_stream_buff_0;
       in_stream_buff_1 <= in_stream_buff_1;
       in_stream_empty <= in_stream_empty;
       in_stream_full <= in_stream_full;
       slice_stream_buff_0 <= slice_stream_buff_0;
       slice_stream_buff_1 <= slice_stream_buff_1;
       slice_stream_empty <= slice_stream_empty;
       slice_stream_full <= slice_stream_full;
       stencil_stream_buff_0 <= stencil_stream_buff_0;
       stencil_stream_buff_1 <= stencil_stream_buff_1;
       stencil_stream_empty <= stencil_stream_empty;
       stencil_stream_full <= stencil_stream_full;
   end
   else if(step) begin
       LB1D_buff <= n38;
       LB1D_in <= n44;
       LB1D_it_1 <= n45;
       LB1D_p_cnt <= n55;
       LB1D_uIn <= n60;
       LB2D_proc_w <= n70;
       LB2D_proc_x <= n77;
       LB2D_proc_y <= n86;
       LB2D_shift_0 <= n91;
       LB2D_shift_1 <= n96;
       LB2D_shift_2 <= n101;
       LB2D_shift_3 <= n106;
       LB2D_shift_4 <= n111;
       LB2D_shift_5 <= n116;
       LB2D_shift_6 <= n121;
       LB2D_shift_7 <= n128;
       LB2D_shift_x <= n134;
       LB2D_shift_y <= n144;
       arg_0_TDATA <= n152;
       arg_0_TVALID <= n159;
       arg_1_TREADY <= n165;
       gb_exit_it_1 <= n173;
       gb_exit_it_2 <= n178;
       gb_exit_it_3 <= n183;
       gb_exit_it_4 <= n188;
       gb_exit_it_5 <= n193;
       gb_exit_it_6 <= n198;
       gb_exit_it_7 <= n203;
       gb_exit_it_8 <= n208;
       gb_p_cnt <= n215;
       gb_pp_it_1 <= n220;
       gb_pp_it_2 <= n225;
       gb_pp_it_3 <= n230;
       gb_pp_it_4 <= n235;
       gb_pp_it_5 <= n240;
       gb_pp_it_6 <= n245;
       gb_pp_it_7 <= n250;
       gb_pp_it_8 <= n255;
       gb_pp_it_9 <= n260;
       in_stream_buff_0 <= n265;
       in_stream_buff_1 <= n270;
       in_stream_empty <= n277;
       in_stream_full <= n284;
       slice_stream_buff_0 <= n371;
       slice_stream_buff_1 <= n377;
       slice_stream_empty <= n384;
       slice_stream_full <= n392;
       stencil_stream_buff_0 <= n560;
       stencil_stream_buff_1 <= n565;
       stencil_stream_empty <= n572;
       stencil_stream_full <= n581;
       LB2D_proc_0 [ LB2D_proc_0_addr0 ] <= LB2D_proc_0_data0;
       LB2D_proc_1 [ LB2D_proc_1_addr0 ] <= LB2D_proc_1_data0;
       LB2D_proc_2 [ LB2D_proc_2_addr0 ] <= LB2D_proc_2_data0;
       LB2D_proc_3 [ LB2D_proc_3_addr0 ] <= LB2D_proc_3_data0;
       LB2D_proc_4 [ LB2D_proc_4_addr0 ] <= LB2D_proc_4_data0;
       LB2D_proc_5 [ LB2D_proc_5_addr0 ] <= LB2D_proc_5_data0;
       LB2D_proc_6 [ LB2D_proc_6_addr0 ] <= LB2D_proc_6_data0;
       LB2D_proc_7 [ LB2D_proc_7_addr0 ] <= LB2D_proc_7_data0;
   end
end
endmodule
