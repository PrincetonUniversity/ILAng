module GB(
arg_0_TREADY,
arg_1_TDATA,
arg_1_TVALID,
LB1D_buff,
LB1D_it_1,
LB1D_p_cnt,
LB2D_proc_w,
LB2D_proc_x,
LB2D_proc_y,
LB2D_shift_0,
LB2D_shift_1,
LB2D_shift_2,
LB2D_shift_3,
LB2D_shift_4,
LB2D_shift_5,
LB2D_shift_6,
LB2D_shift_7,
LB2D_shift_x,
LB2D_shift_y,
arg_0_TDATA,
arg_0_TVALID,
arg_1_TREADY,
gb_exit_it_1,
gb_exit_it_2,
gb_exit_it_3,
gb_exit_it_4,
gb_exit_it_5,
gb_exit_it_6,
gb_exit_it_7,
gb_exit_it_8,
gb_p_cnt,
gb_pp_it_1,
gb_pp_it_2,
gb_pp_it_3,
gb_pp_it_4,
gb_pp_it_5,
gb_pp_it_6,
gb_pp_it_7,
gb_pp_it_8,
gb_pp_it_9,
in_stream_buff_0,
in_stream_buff_1,
in_stream_empty,
in_stream_full,
slice_stream_buff_0,
slice_stream_buff_1,
slice_stream_empty,
slice_stream_full,
stencil_stream_buff_0,
stencil_stream_buff_1,
stencil_stream_empty,
stencil_stream_full,
clk,rst,
step
);
input            arg_0_TREADY;
input      [7:0] arg_1_TDATA;
input            arg_1_TVALID;
input clk;
input rst;
input step;
output      [7:0] LB1D_buff;
output            LB1D_it_1;
output     [18:0] LB1D_p_cnt;
output     [63:0] LB2D_proc_w;
output      [8:0] LB2D_proc_x;
output      [9:0] LB2D_proc_y;
output     [71:0] LB2D_shift_0;
output     [71:0] LB2D_shift_1;
output     [71:0] LB2D_shift_2;
output     [71:0] LB2D_shift_3;
output     [71:0] LB2D_shift_4;
output     [71:0] LB2D_shift_5;
output     [71:0] LB2D_shift_6;
output     [71:0] LB2D_shift_7;
output      [8:0] LB2D_shift_x;
output      [9:0] LB2D_shift_y;
output      [7:0] arg_0_TDATA;
output            arg_0_TVALID;
output            arg_1_TREADY;
output            gb_exit_it_1;
output            gb_exit_it_2;
output            gb_exit_it_3;
output            gb_exit_it_4;
output            gb_exit_it_5;
output            gb_exit_it_6;
output            gb_exit_it_7;
output            gb_exit_it_8;
output     [18:0] gb_p_cnt;
output            gb_pp_it_1;
output            gb_pp_it_2;
output            gb_pp_it_3;
output            gb_pp_it_4;
output            gb_pp_it_5;
output            gb_pp_it_6;
output            gb_pp_it_7;
output            gb_pp_it_8;
output            gb_pp_it_9;
output      [7:0] in_stream_buff_0;
output      [7:0] in_stream_buff_1;
output            in_stream_empty;
output            in_stream_full;
output     [71:0] slice_stream_buff_0;
output     [71:0] slice_stream_buff_1;
output            slice_stream_empty;
output            slice_stream_full;
output    [647:0] stencil_stream_buff_0;
output    [647:0] stencil_stream_buff_1;
output            stencil_stream_empty;
output            stencil_stream_full;
reg      [7:0] LB1D_buff;
reg            LB1D_it_1;
reg     [18:0] LB1D_p_cnt;
reg     [63:0] LB2D_proc_w;
reg      [8:0] LB2D_proc_x;
reg      [9:0] LB2D_proc_y;
reg     [71:0] LB2D_shift_0;
reg     [71:0] LB2D_shift_1;
reg     [71:0] LB2D_shift_2;
reg     [71:0] LB2D_shift_3;
reg     [71:0] LB2D_shift_4;
reg     [71:0] LB2D_shift_5;
reg     [71:0] LB2D_shift_6;
reg     [71:0] LB2D_shift_7;
reg      [8:0] LB2D_shift_x;
reg      [9:0] LB2D_shift_y;
reg      [7:0] arg_0_TDATA;
reg            arg_0_TVALID;
reg            arg_1_TREADY;
reg            gb_exit_it_1;
reg            gb_exit_it_2;
reg            gb_exit_it_3;
reg            gb_exit_it_4;
reg            gb_exit_it_5;
reg            gb_exit_it_6;
reg            gb_exit_it_7;
reg            gb_exit_it_8;
reg     [18:0] gb_p_cnt;
reg            gb_pp_it_1;
reg            gb_pp_it_2;
reg            gb_pp_it_3;
reg            gb_pp_it_4;
reg            gb_pp_it_5;
reg            gb_pp_it_6;
reg            gb_pp_it_7;
reg            gb_pp_it_8;
reg            gb_pp_it_9;
reg      [7:0] in_stream_buff_0;
reg      [7:0] in_stream_buff_1;
reg            in_stream_empty;
reg            in_stream_full;
reg     [71:0] slice_stream_buff_0;
reg     [71:0] slice_stream_buff_1;
reg            slice_stream_empty;
reg            slice_stream_full;
reg    [647:0] stencil_stream_buff_0;
reg    [647:0] stencil_stream_buff_1;
reg            stencil_stream_empty;
reg            stencil_stream_full;
wire            arg_0_TREADY;
wire      [7:0] arg_1_TDATA;
wire            arg_1_TVALID;
wire            n0;
wire            n1;
wire            n2;
wire            n3;
wire            n4;
wire            n5;
wire            n6;
wire            n7;
wire            n8;
wire            n9;
wire            n10;
wire            n11;
wire            n12;
wire            n13;
wire            n14;
wire            n15;
wire            n16;
wire            n17;
wire            n18;
wire            n19;
wire            n20;
wire            n21;
wire            n22;
wire            n23;
wire            n24;
wire            n25;
wire            n26;
wire            n27;
wire            n28;
wire            n29;
wire            n30;
wire            n31;
wire            n32;
wire            n33;
wire            n34;
wire            n35;
wire            n36;
wire            n37;
wire      [7:0] n38;
wire      [7:0] n39;
wire      [7:0] n40;
wire      [7:0] n41;
wire      [7:0] n42;
wire      [7:0] n43;
wire            n44;
wire            n45;
wire            n46;
wire     [18:0] n47;
wire     [18:0] n48;
wire            n49;
wire     [18:0] n50;
wire     [18:0] n51;
wire     [18:0] n52;
wire     [18:0] n53;
wire     [18:0] n54;
wire     [18:0] n55;
wire     [18:0] n56;
wire     [18:0] n57;
wire            n58;
wire            n59;
wire     [63:0] n60;
wire     [63:0] n61;
wire     [63:0] n62;
wire     [63:0] n63;
wire     [63:0] n64;
wire     [63:0] n65;
wire     [63:0] n66;
wire     [63:0] n67;
wire     [63:0] n68;
wire            n69;
wire            n70;
wire            n71;
wire      [8:0] n72;
wire      [8:0] n73;
wire      [8:0] n74;
wire      [8:0] n75;
wire      [8:0] n76;
wire      [8:0] n77;
wire      [8:0] n78;
wire      [8:0] n79;
wire            n80;
wire      [9:0] n81;
wire      [9:0] n82;
wire      [9:0] n83;
wire      [9:0] n84;
wire      [9:0] n85;
wire      [9:0] n86;
wire      [9:0] n87;
wire            n88;
wire     [71:0] n89;
wire     [71:0] n90;
wire     [71:0] n91;
wire     [71:0] n92;
wire     [71:0] n93;
wire     [71:0] n94;
wire     [71:0] n95;
wire     [71:0] n96;
wire     [71:0] n97;
wire     [71:0] n98;
wire     [71:0] n99;
wire     [71:0] n100;
wire     [71:0] n101;
wire     [71:0] n102;
wire     [71:0] n103;
wire     [71:0] n104;
wire     [71:0] n105;
wire     [71:0] n106;
wire     [71:0] n107;
wire     [71:0] n108;
wire     [71:0] n109;
wire     [71:0] n110;
wire     [71:0] n111;
wire     [71:0] n112;
wire     [71:0] n113;
wire     [71:0] n114;
wire     [71:0] n115;
wire     [71:0] n116;
wire     [71:0] n117;
wire     [71:0] n118;
wire     [71:0] n119;
wire     [71:0] n120;
wire     [71:0] n121;
wire     [71:0] n122;
wire     [71:0] n123;
wire     [71:0] n124;
wire     [71:0] n125;
wire     [71:0] n126;
wire     [71:0] n127;
wire     [71:0] n128;
wire     [71:0] n129;
wire     [71:0] n130;
wire     [71:0] n131;
wire     [71:0] n132;
wire     [71:0] n133;
wire     [71:0] n134;
wire     [71:0] n135;
wire     [71:0] n136;
wire     [71:0] n137;
wire      [8:0] n138;
wire      [8:0] n139;
wire      [8:0] n140;
wire      [8:0] n141;
wire      [8:0] n142;
wire      [8:0] n143;
wire      [8:0] n144;
wire            n145;
wire            n146;
wire      [9:0] n147;
wire      [9:0] n148;
wire      [9:0] n149;
wire      [9:0] n150;
wire      [9:0] n151;
wire      [9:0] n152;
wire      [9:0] n153;
wire      [9:0] n154;
wire      [9:0] n155;
wire            n156;
wire    [647:0] n157;
wire      [7:0] n158;
wire      [7:0] n159;
wire      [7:0] n160;
wire      [7:0] n161;
wire      [7:0] n162;
wire      [7:0] n163;
wire      [7:0] n164;
wire            n165;
wire            n166;
wire            n167;
wire            n168;
wire            n169;
wire            n170;
wire            n171;
wire            n172;
wire            n173;
wire            n174;
wire            n175;
wire            n176;
wire            n177;
wire            n178;
wire            n179;
wire     [18:0] n180;
wire            n181;
wire            n182;
wire            n183;
wire            n184;
wire            n185;
wire            n186;
wire            n187;
wire            n188;
wire            n189;
wire            n190;
wire            n191;
wire            n192;
wire            n193;
wire            n194;
wire            n195;
wire            n196;
wire            n197;
wire            n198;
wire            n199;
wire            n200;
wire            n201;
wire            n202;
wire            n203;
wire            n204;
wire            n205;
wire            n206;
wire            n207;
wire            n208;
wire            n209;
wire            n210;
wire            n211;
wire            n212;
wire            n213;
wire            n214;
wire            n215;
wire            n216;
wire            n217;
wire            n218;
wire            n219;
wire            n220;
wire            n221;
wire            n222;
wire            n223;
wire            n224;
wire            n225;
wire            n226;
wire            n227;
wire            n228;
wire            n229;
wire            n230;
wire            n231;
wire     [18:0] n232;
wire     [18:0] n233;
wire     [18:0] n234;
wire     [18:0] n235;
wire     [18:0] n236;
wire     [18:0] n237;
wire     [18:0] n238;
wire            n239;
wire            n240;
wire            n241;
wire            n242;
wire            n243;
wire            n244;
wire            n245;
wire            n246;
wire            n247;
wire            n248;
wire            n249;
wire            n250;
wire            n251;
wire            n252;
wire            n253;
wire            n254;
wire            n255;
wire            n256;
wire            n257;
wire            n258;
wire            n259;
wire            n260;
wire            n261;
wire            n262;
wire            n263;
wire            n264;
wire            n265;
wire            n266;
wire            n267;
wire            n268;
wire            n269;
wire            n270;
wire            n271;
wire            n272;
wire            n273;
wire            n274;
wire            n275;
wire            n276;
wire            n277;
wire            n278;
wire            n279;
wire            n280;
wire            n281;
wire            n282;
wire            n283;
wire            n284;
wire            n285;
wire            n286;
wire            n287;
wire            n288;
wire            n289;
wire            n290;
wire            n291;
wire            n292;
wire      [7:0] n293;
wire      [7:0] n294;
wire      [7:0] n295;
wire      [7:0] n296;
wire      [7:0] n297;
wire      [7:0] n298;
wire      [7:0] n299;
wire      [7:0] n300;
wire      [7:0] n301;
wire      [7:0] n302;
wire      [7:0] n303;
wire      [7:0] n304;
wire            n305;
wire            n306;
wire            n307;
wire            n308;
wire            n309;
wire            n310;
wire            n311;
wire            n312;
wire            n313;
wire            n314;
wire            n315;
wire            n316;
wire            n317;
wire            n318;
wire            n319;
wire            n320;
wire      [7:0] n321;
wire            n322;
wire      [7:0] n323;
wire            n324;
wire      [7:0] n325;
wire            n326;
wire      [7:0] n327;
wire            n328;
wire      [7:0] n329;
wire            n330;
wire      [7:0] n331;
wire            n332;
wire      [7:0] n333;
wire            n334;
wire      [7:0] n335;
wire      [7:0] n336;
wire      [7:0] n337;
wire      [7:0] n338;
wire      [7:0] n339;
wire      [7:0] n340;
wire      [7:0] n341;
wire      [7:0] n342;
wire      [7:0] n343;
wire      [7:0] n344;
wire      [7:0] n345;
wire      [7:0] n346;
wire      [7:0] n347;
wire      [7:0] n348;
wire      [7:0] n349;
wire      [7:0] n350;
wire      [7:0] n351;
wire      [7:0] n352;
wire      [7:0] n353;
wire      [7:0] n354;
wire      [7:0] n355;
wire      [7:0] n356;
wire      [7:0] n357;
wire      [7:0] n358;
wire      [7:0] n359;
wire      [7:0] n360;
wire      [7:0] n361;
wire      [7:0] n362;
wire      [7:0] n363;
wire      [7:0] n364;
wire      [7:0] n365;
wire      [7:0] n366;
wire      [7:0] n367;
wire      [7:0] n368;
wire      [7:0] n369;
wire      [7:0] n370;
wire      [7:0] n371;
wire      [7:0] n372;
wire      [7:0] n373;
wire      [7:0] n374;
wire      [7:0] n375;
wire      [7:0] n376;
wire      [7:0] n377;
wire      [7:0] n378;
wire      [7:0] n379;
wire      [7:0] n380;
wire      [7:0] n381;
wire      [7:0] n382;
wire      [7:0] n383;
wire      [7:0] n384;
wire      [7:0] n385;
wire      [7:0] n386;
wire      [7:0] n387;
wire      [7:0] n388;
wire      [7:0] n389;
wire      [7:0] n390;
wire      [7:0] n391;
wire      [7:0] n392;
wire     [15:0] n393;
wire     [23:0] n394;
wire     [31:0] n395;
wire     [39:0] n396;
wire     [47:0] n397;
wire     [55:0] n398;
wire     [63:0] n399;
wire     [71:0] n400;
wire     [71:0] n401;
wire     [71:0] n402;
wire     [71:0] n403;
wire     [71:0] n404;
wire     [71:0] n405;
wire     [71:0] n406;
wire     [71:0] n407;
wire     [71:0] n408;
wire     [71:0] n409;
wire     [71:0] n410;
wire     [71:0] n411;
wire     [71:0] n412;
wire     [71:0] n413;
wire     [71:0] n414;
wire            n415;
wire            n416;
wire            n417;
wire            n418;
wire            n419;
wire            n420;
wire            n421;
wire            n422;
wire            n423;
wire            n424;
wire            n425;
wire            n426;
wire            n427;
wire            n428;
wire            n429;
wire            n430;
wire            n431;
wire            n432;
wire      [7:0] n433;
wire      [7:0] n434;
wire      [7:0] n435;
wire      [7:0] n436;
wire      [7:0] n437;
wire      [7:0] n438;
wire      [7:0] n439;
wire      [7:0] n440;
wire      [7:0] n441;
wire     [15:0] n442;
wire     [23:0] n443;
wire     [31:0] n444;
wire     [39:0] n445;
wire     [47:0] n446;
wire     [55:0] n447;
wire     [63:0] n448;
wire     [71:0] n449;
wire      [7:0] n450;
wire      [7:0] n451;
wire      [7:0] n452;
wire      [7:0] n453;
wire      [7:0] n454;
wire      [7:0] n455;
wire      [7:0] n456;
wire      [7:0] n457;
wire      [7:0] n458;
wire     [15:0] n459;
wire     [23:0] n460;
wire     [31:0] n461;
wire     [39:0] n462;
wire     [47:0] n463;
wire     [55:0] n464;
wire     [63:0] n465;
wire     [71:0] n466;
wire      [7:0] n467;
wire      [7:0] n468;
wire      [7:0] n469;
wire      [7:0] n470;
wire      [7:0] n471;
wire      [7:0] n472;
wire      [7:0] n473;
wire      [7:0] n474;
wire      [7:0] n475;
wire     [15:0] n476;
wire     [23:0] n477;
wire     [31:0] n478;
wire     [39:0] n479;
wire     [47:0] n480;
wire     [55:0] n481;
wire     [63:0] n482;
wire     [71:0] n483;
wire      [7:0] n484;
wire      [7:0] n485;
wire      [7:0] n486;
wire      [7:0] n487;
wire      [7:0] n488;
wire      [7:0] n489;
wire      [7:0] n490;
wire      [7:0] n491;
wire      [7:0] n492;
wire     [15:0] n493;
wire     [23:0] n494;
wire     [31:0] n495;
wire     [39:0] n496;
wire     [47:0] n497;
wire     [55:0] n498;
wire     [63:0] n499;
wire     [71:0] n500;
wire      [7:0] n501;
wire      [7:0] n502;
wire      [7:0] n503;
wire      [7:0] n504;
wire      [7:0] n505;
wire      [7:0] n506;
wire      [7:0] n507;
wire      [7:0] n508;
wire      [7:0] n509;
wire     [15:0] n510;
wire     [23:0] n511;
wire     [31:0] n512;
wire     [39:0] n513;
wire     [47:0] n514;
wire     [55:0] n515;
wire     [63:0] n516;
wire     [71:0] n517;
wire      [7:0] n518;
wire      [7:0] n519;
wire      [7:0] n520;
wire      [7:0] n521;
wire      [7:0] n522;
wire      [7:0] n523;
wire      [7:0] n524;
wire      [7:0] n525;
wire      [7:0] n526;
wire     [15:0] n527;
wire     [23:0] n528;
wire     [31:0] n529;
wire     [39:0] n530;
wire     [47:0] n531;
wire     [55:0] n532;
wire     [63:0] n533;
wire     [71:0] n534;
wire      [7:0] n535;
wire      [7:0] n536;
wire      [7:0] n537;
wire      [7:0] n538;
wire      [7:0] n539;
wire      [7:0] n540;
wire      [7:0] n541;
wire      [7:0] n542;
wire      [7:0] n543;
wire     [15:0] n544;
wire     [23:0] n545;
wire     [31:0] n546;
wire     [39:0] n547;
wire     [47:0] n548;
wire     [55:0] n549;
wire     [63:0] n550;
wire     [71:0] n551;
wire      [7:0] n552;
wire      [7:0] n553;
wire      [7:0] n554;
wire      [7:0] n555;
wire      [7:0] n556;
wire      [7:0] n557;
wire      [7:0] n558;
wire      [7:0] n559;
wire      [7:0] n560;
wire     [15:0] n561;
wire     [23:0] n562;
wire     [31:0] n563;
wire     [39:0] n564;
wire     [47:0] n565;
wire     [55:0] n566;
wire     [63:0] n567;
wire     [71:0] n568;
wire      [7:0] n569;
wire      [7:0] n570;
wire      [7:0] n571;
wire      [7:0] n572;
wire      [7:0] n573;
wire      [7:0] n574;
wire      [7:0] n575;
wire      [7:0] n576;
wire      [7:0] n577;
wire     [15:0] n578;
wire     [23:0] n579;
wire     [31:0] n580;
wire     [39:0] n581;
wire     [47:0] n582;
wire     [55:0] n583;
wire     [63:0] n584;
wire     [71:0] n585;
wire    [143:0] n586;
wire    [215:0] n587;
wire    [287:0] n588;
wire    [359:0] n589;
wire    [431:0] n590;
wire    [503:0] n591;
wire    [575:0] n592;
wire    [647:0] n593;
wire    [647:0] n594;
wire    [647:0] n595;
wire    [647:0] n596;
wire    [647:0] n597;
wire    [647:0] n598;
wire    [647:0] n599;
wire    [647:0] n600;
wire    [647:0] n601;
wire    [647:0] n602;
wire    [647:0] n603;
wire    [647:0] n604;
wire    [647:0] n605;
wire    [647:0] n606;
wire            n607;
wire            n608;
wire            n609;
wire            n610;
wire            n611;
wire            n612;
wire            n613;
wire            n614;
wire            n615;
wire            n616;
wire            n617;
wire            n618;
wire            n619;
wire            n620;
wire            n621;
wire            n622;
wire            n623;
wire            n624;
wire      [8:0] LB2D_proc_0_addr0;
wire      [7:0] LB2D_proc_0_data0;
wire            n625;
wire            n626;
wire            n627;
wire            n628;
wire            n629;
wire            n630;
wire            n631;
wire            n632;
wire            n633;
wire            n634;
wire            n635;
wire            n636;
wire            n637;
wire            n638;
wire            n639;
wire            n640;
wire            n641;
wire            n642;
wire            n643;
wire      [8:0] LB2D_proc_1_addr0;
wire      [7:0] LB2D_proc_1_data0;
wire            n644;
wire            n645;
wire            n646;
wire      [8:0] LB2D_proc_2_addr0;
wire      [7:0] LB2D_proc_2_data0;
wire            n647;
wire            n648;
wire            n649;
wire      [8:0] LB2D_proc_3_addr0;
wire      [7:0] LB2D_proc_3_data0;
wire            n650;
wire            n651;
wire            n652;
wire      [8:0] LB2D_proc_4_addr0;
wire      [7:0] LB2D_proc_4_data0;
wire            n653;
wire            n654;
wire            n655;
wire      [8:0] LB2D_proc_5_addr0;
wire      [7:0] LB2D_proc_5_data0;
wire            n656;
wire            n657;
wire            n658;
wire      [8:0] LB2D_proc_6_addr0;
wire      [7:0] LB2D_proc_6_data0;
wire            n659;
wire            n660;
wire            n661;
wire      [8:0] LB2D_proc_7_addr0;
wire      [7:0] LB2D_proc_7_data0;
wire            n662;
wire            n663;
wire            n664;
wire            n665;
reg      [7:0] LB2D_proc_0[511:0];
reg      [7:0] LB2D_proc_1[511:0];
reg      [7:0] LB2D_proc_2[511:0];
reg      [7:0] LB2D_proc_3[511:0];
reg      [7:0] LB2D_proc_4[511:0];
reg      [7:0] LB2D_proc_5[511:0];
reg      [7:0] LB2D_proc_6[511:0];
reg      [7:0] LB2D_proc_7[511:0];
wire clk;
wire rst;
wire step;
assign n0 =  ( arg_0_TREADY ) == ( 1'd1 )  ;
assign n1 =  ( arg_0_TVALID ) == ( 1'd1 )  ;
assign n2 =  ( n0 ) & ( n1 )  ;
assign n3 =  ( arg_1_TVALID ) == ( 1'd0 )  ;
assign n4 =  ( n2 ) & ( n3 )  ;
assign n5 =  ( arg_1_TREADY ) == ( 1'd1 )  ;
assign n6 =  ( arg_1_TVALID ) == ( 1'd1 )  ;
assign n7 =  ( n5 ) & ( n6 )  ;
assign n8 =  ( arg_0_TREADY ) == ( 1'd0 )  ;
assign n9 =  ( n7 ) & ( n8 )  ;
assign n10 =  ( arg_0_TVALID ) == ( 1'd0 )  ;
assign n11 =  ( gb_exit_it_1 ) == ( 1'd0 )  ;
assign n12 =  ( stencil_stream_empty ) == ( 1'd0 )  ;
assign n13 =  ( n11 ) & ( n12 )  ;
assign n14 =  ( gb_exit_it_1 ) == ( 1'd1 )  ;
assign n15 =  ( gb_exit_it_8 ) == ( 1'd0 )  ;
assign n16 =  ( n14 ) & ( n15 )  ;
assign n17 =  ( n13 ) | ( n16 )  ;
assign n18 =  ( n10 ) & ( n17 )  ;
assign n19 =  ( slice_stream_empty ) == ( 1'd0 )  ;
assign n20 =  ( LB2D_shift_x ) != ( 9'd488 )  ;
assign n21 =  ( n19 ) & ( n20 )  ;
assign n22 =  ( stencil_stream_full ) == ( 1'd0 )  ;
assign n23 =  ( LB2D_shift_x ) < ( 9'd8 )  ;
assign n24 =  ( n22 ) | ( n23 )  ;
assign n25 =  ( n21 ) & ( n24 )  ;
assign n26 =  ( in_stream_empty ) == ( 1'd0 )  ;
assign n27 =  ( LB2D_proc_x ) != ( 9'd488 )  ;
assign n28 =  ( n26 ) & ( n27 )  ;
assign n29 =  ( slice_stream_full ) == ( 1'd0 )  ;
assign n30 =  ( LB2D_proc_y ) < ( 10'd8 )  ;
assign n31 =  ( n29 ) | ( n30 )  ;
assign n32 =  ( n28 ) & ( n31 )  ;
assign n33 =  ( arg_1_TREADY ) == ( 1'd0 )  ;
assign n34 =  ( in_stream_full ) == ( 1'd0 )  ;
assign n35 =  ( n33 ) & ( n34 )  ;
assign n36 =  ( LB1D_it_1 ) == ( 1'd1 )  ;
assign n37 =  ( n35 ) & ( n36 )  ;
assign n38 =  ( n37 ) ? ( LB1D_buff ) : ( LB1D_buff ) ;
assign n39 =  ( n32 ) ? ( LB1D_buff ) : ( n38 ) ;
assign n40 =  ( n25 ) ? ( LB1D_buff ) : ( n39 ) ;
assign n41 =  ( n18 ) ? ( LB1D_buff ) : ( n40 ) ;
assign n42 =  ( n9 ) ? ( arg_1_TDATA ) : ( n41 ) ;
assign n43 =  ( n4 ) ? ( arg_1_TDATA ) : ( n42 ) ;
assign n44 =  ( LB1D_it_1 ) == ( 1'd0 )  ;
assign n45 =  ( n35 ) & ( n44 )  ;
assign n46 =  ( n45 ) ? ( 1'd1 ) : ( LB1D_it_1 ) ;
assign n47 =  ( LB1D_p_cnt ) + ( 19'd1 )  ;
assign n48 =  ( 19'd316224 ) - ( 19'd1 )  ;
assign n49 =  ( LB1D_p_cnt ) == ( n48 )  ;
assign n50 =  ( n49 ) ? ( 19'd0 ) : ( n47 ) ;
assign n51 =  ( n37 ) ? ( n50 ) : ( LB1D_p_cnt ) ;
assign n52 =  ( n45 ) ? ( n47 ) : ( n51 ) ;
assign n53 =  ( n32 ) ? ( LB1D_p_cnt ) : ( n52 ) ;
assign n54 =  ( n25 ) ? ( LB1D_p_cnt ) : ( n53 ) ;
assign n55 =  ( n18 ) ? ( LB1D_p_cnt ) : ( n54 ) ;
assign n56 =  ( n9 ) ? ( LB1D_p_cnt ) : ( n55 ) ;
assign n57 =  ( n4 ) ? ( LB1D_p_cnt ) : ( n56 ) ;
assign n58 =  ( LB2D_proc_w ) < ( 64'd7 )  ;
assign n59 =  ( LB2D_proc_x ) < ( 9'd488 )  ;
assign n60 =  ( LB2D_proc_w ) + ( 64'd1 )  ;
assign n61 =  ( n59 ) ? ( LB2D_proc_w ) : ( n60 ) ;
assign n62 =  ( n58 ) ? ( n61 ) : ( 64'd0 ) ;
assign n63 =  ( n37 ) ? ( LB2D_proc_w ) : ( LB2D_proc_w ) ;
assign n64 =  ( n32 ) ? ( n62 ) : ( n63 ) ;
assign n65 =  ( n25 ) ? ( LB2D_proc_w ) : ( n64 ) ;
assign n66 =  ( n18 ) ? ( LB2D_proc_w ) : ( n65 ) ;
assign n67 =  ( n9 ) ? ( LB2D_proc_w ) : ( n66 ) ;
assign n68 =  ( n4 ) ? ( LB2D_proc_w ) : ( n67 ) ;
assign n69 =  ( LB2D_proc_x ) == ( 9'd488 )  ;
assign n70 =  ( n26 ) & ( n69 )  ;
assign n71 =  ( n70 ) & ( n31 )  ;
assign n72 =  ( LB2D_proc_x ) + ( 9'd1 )  ;
assign n73 =  ( n37 ) ? ( LB2D_proc_x ) : ( LB2D_proc_x ) ;
assign n74 =  ( n32 ) ? ( n72 ) : ( n73 ) ;
assign n75 =  ( n71 ) ? ( 9'd0 ) : ( n74 ) ;
assign n76 =  ( n25 ) ? ( LB2D_proc_x ) : ( n75 ) ;
assign n77 =  ( n18 ) ? ( LB2D_proc_x ) : ( n76 ) ;
assign n78 =  ( n9 ) ? ( LB2D_proc_x ) : ( n77 ) ;
assign n79 =  ( n4 ) ? ( LB2D_proc_x ) : ( n78 ) ;
assign n80 =  ( LB2D_proc_y ) < ( 10'd488 )  ;
assign n81 =  ( n80 ) ? ( LB2D_proc_y ) : ( 10'd488 ) ;
assign n82 =  ( n37 ) ? ( LB2D_proc_y ) : ( LB2D_proc_y ) ;
assign n83 =  ( n32 ) ? ( n81 ) : ( n82 ) ;
assign n84 =  ( n25 ) ? ( LB2D_proc_y ) : ( n83 ) ;
assign n85 =  ( n18 ) ? ( LB2D_proc_y ) : ( n84 ) ;
assign n86 =  ( n9 ) ? ( LB2D_proc_y ) : ( n85 ) ;
assign n87 =  ( n4 ) ? ( LB2D_proc_y ) : ( n86 ) ;
assign n88 =  ( slice_stream_full ) == ( 1'd1 )  ;
assign n89 =  ( n88 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n90 =  ( n37 ) ? ( LB2D_shift_0 ) : ( LB2D_shift_0 ) ;
assign n91 =  ( n32 ) ? ( LB2D_shift_0 ) : ( n90 ) ;
assign n92 =  ( n25 ) ? ( n89 ) : ( n91 ) ;
assign n93 =  ( n18 ) ? ( LB2D_shift_0 ) : ( n92 ) ;
assign n94 =  ( n9 ) ? ( LB2D_shift_0 ) : ( n93 ) ;
assign n95 =  ( n4 ) ? ( LB2D_shift_0 ) : ( n94 ) ;
assign n96 =  ( n37 ) ? ( LB2D_shift_1 ) : ( LB2D_shift_1 ) ;
assign n97 =  ( n32 ) ? ( LB2D_shift_1 ) : ( n96 ) ;
assign n98 =  ( n25 ) ? ( LB2D_shift_0 ) : ( n97 ) ;
assign n99 =  ( n18 ) ? ( LB2D_shift_1 ) : ( n98 ) ;
assign n100 =  ( n9 ) ? ( LB2D_shift_1 ) : ( n99 ) ;
assign n101 =  ( n4 ) ? ( LB2D_shift_1 ) : ( n100 ) ;
assign n102 =  ( n37 ) ? ( LB2D_shift_2 ) : ( LB2D_shift_2 ) ;
assign n103 =  ( n32 ) ? ( LB2D_shift_2 ) : ( n102 ) ;
assign n104 =  ( n25 ) ? ( LB2D_shift_1 ) : ( n103 ) ;
assign n105 =  ( n18 ) ? ( LB2D_shift_2 ) : ( n104 ) ;
assign n106 =  ( n9 ) ? ( LB2D_shift_2 ) : ( n105 ) ;
assign n107 =  ( n4 ) ? ( LB2D_shift_2 ) : ( n106 ) ;
assign n108 =  ( n37 ) ? ( LB2D_shift_3 ) : ( LB2D_shift_3 ) ;
assign n109 =  ( n32 ) ? ( LB2D_shift_3 ) : ( n108 ) ;
assign n110 =  ( n25 ) ? ( LB2D_shift_2 ) : ( n109 ) ;
assign n111 =  ( n18 ) ? ( LB2D_shift_3 ) : ( n110 ) ;
assign n112 =  ( n9 ) ? ( LB2D_shift_3 ) : ( n111 ) ;
assign n113 =  ( n4 ) ? ( LB2D_shift_3 ) : ( n112 ) ;
assign n114 =  ( n37 ) ? ( LB2D_shift_4 ) : ( LB2D_shift_4 ) ;
assign n115 =  ( n32 ) ? ( LB2D_shift_4 ) : ( n114 ) ;
assign n116 =  ( n25 ) ? ( LB2D_shift_3 ) : ( n115 ) ;
assign n117 =  ( n18 ) ? ( LB2D_shift_4 ) : ( n116 ) ;
assign n118 =  ( n9 ) ? ( LB2D_shift_4 ) : ( n117 ) ;
assign n119 =  ( n4 ) ? ( LB2D_shift_4 ) : ( n118 ) ;
assign n120 =  ( n37 ) ? ( LB2D_shift_5 ) : ( LB2D_shift_5 ) ;
assign n121 =  ( n32 ) ? ( LB2D_shift_5 ) : ( n120 ) ;
assign n122 =  ( n25 ) ? ( LB2D_shift_4 ) : ( n121 ) ;
assign n123 =  ( n18 ) ? ( LB2D_shift_5 ) : ( n122 ) ;
assign n124 =  ( n9 ) ? ( LB2D_shift_5 ) : ( n123 ) ;
assign n125 =  ( n4 ) ? ( LB2D_shift_5 ) : ( n124 ) ;
assign n126 =  ( n37 ) ? ( LB2D_shift_6 ) : ( LB2D_shift_6 ) ;
assign n127 =  ( n32 ) ? ( LB2D_shift_6 ) : ( n126 ) ;
assign n128 =  ( n25 ) ? ( LB2D_shift_5 ) : ( n127 ) ;
assign n129 =  ( n18 ) ? ( LB2D_shift_6 ) : ( n128 ) ;
assign n130 =  ( n9 ) ? ( LB2D_shift_6 ) : ( n129 ) ;
assign n131 =  ( n4 ) ? ( LB2D_shift_6 ) : ( n130 ) ;
assign n132 =  ( n37 ) ? ( LB2D_shift_7 ) : ( LB2D_shift_7 ) ;
assign n133 =  ( n32 ) ? ( LB2D_shift_7 ) : ( n132 ) ;
assign n134 =  ( n25 ) ? ( LB2D_shift_6 ) : ( n133 ) ;
assign n135 =  ( n18 ) ? ( LB2D_shift_7 ) : ( n134 ) ;
assign n136 =  ( n9 ) ? ( LB2D_shift_7 ) : ( n135 ) ;
assign n137 =  ( n4 ) ? ( LB2D_shift_7 ) : ( n136 ) ;
assign n138 =  ( LB2D_shift_x ) + ( 9'd1 )  ;
assign n139 =  ( n37 ) ? ( LB2D_shift_x ) : ( LB2D_shift_x ) ;
assign n140 =  ( n32 ) ? ( LB2D_shift_x ) : ( n139 ) ;
assign n141 =  ( n25 ) ? ( n138 ) : ( n140 ) ;
assign n142 =  ( n18 ) ? ( LB2D_shift_x ) : ( n141 ) ;
assign n143 =  ( n9 ) ? ( LB2D_shift_x ) : ( n142 ) ;
assign n144 =  ( n4 ) ? ( LB2D_shift_x ) : ( n143 ) ;
assign n145 =  ( LB2D_shift_y ) < ( 10'd480 )  ;
assign n146 =  ( LB2D_shift_x ) < ( 9'd488 )  ;
assign n147 =  ( LB2D_shift_y ) + ( 10'd1 )  ;
assign n148 =  ( n146 ) ? ( LB2D_shift_y ) : ( n147 ) ;
assign n149 =  ( n145 ) ? ( n148 ) : ( 10'd480 ) ;
assign n150 =  ( n37 ) ? ( LB2D_shift_y ) : ( LB2D_shift_y ) ;
assign n151 =  ( n32 ) ? ( LB2D_shift_y ) : ( n150 ) ;
assign n152 =  ( n25 ) ? ( n149 ) : ( n151 ) ;
assign n153 =  ( n18 ) ? ( LB2D_shift_y ) : ( n152 ) ;
assign n154 =  ( n9 ) ? ( LB2D_shift_y ) : ( n153 ) ;
assign n155 =  ( n4 ) ? ( LB2D_shift_y ) : ( n154 ) ;
assign n156 =  ( stencil_stream_full ) == ( 1'd1 )  ;
assign n157 =  ( n156 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_0 ) ;
//assign n158 = gb_fun(n157) ;
gb_fun gb_fun_U (
        .stencil (n157),
        .result (n158)
        );

assign n159 =  ( n37 ) ? ( arg_0_TDATA ) : ( arg_0_TDATA ) ;
assign n160 =  ( n32 ) ? ( arg_0_TDATA ) : ( n159 ) ;
assign n161 =  ( n25 ) ? ( arg_0_TDATA ) : ( n160 ) ;
assign n162 =  ( n18 ) ? ( n158 ) : ( n161 ) ;
assign n163 =  ( n9 ) ? ( arg_0_TDATA ) : ( n162 ) ;
assign n164 =  ( n4 ) ? ( arg_0_TDATA ) : ( n163 ) ;
assign n165 =  ( gb_pp_it_8 ) == ( 1'd1 )  ;
assign n166 =  ( n165 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n167 =  ( n37 ) ? ( arg_0_TVALID ) : ( arg_0_TVALID ) ;
assign n168 =  ( n32 ) ? ( arg_0_TVALID ) : ( n167 ) ;
assign n169 =  ( n25 ) ? ( arg_0_TVALID ) : ( n168 ) ;
assign n170 =  ( n18 ) ? ( n166 ) : ( n169 ) ;
assign n171 =  ( n9 ) ? ( arg_0_TVALID ) : ( n170 ) ;
assign n172 =  ( n4 ) ? ( 1'd0 ) : ( n171 ) ;
assign n173 =  ( n37 ) ? ( 1'd1 ) : ( arg_1_TREADY ) ;
assign n174 =  ( n45 ) ? ( 1'd1 ) : ( n173 ) ;
assign n175 =  ( n32 ) ? ( arg_1_TREADY ) : ( n174 ) ;
assign n176 =  ( n25 ) ? ( arg_1_TREADY ) : ( n175 ) ;
assign n177 =  ( n18 ) ? ( arg_1_TREADY ) : ( n176 ) ;
assign n178 =  ( n9 ) ? ( 1'd0 ) : ( n177 ) ;
assign n179 =  ( n4 ) ? ( 1'd0 ) : ( n178 ) ;
assign n180 =  ( gb_p_cnt ) + ( 19'd1 )  ;
assign n181 =  ( n180 ) == ( 19'd307200 )  ;
assign n182 =  ( n181 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n183 =  ( n37 ) ? ( gb_exit_it_1 ) : ( gb_exit_it_1 ) ;
assign n184 =  ( n32 ) ? ( gb_exit_it_1 ) : ( n183 ) ;
assign n185 =  ( n25 ) ? ( gb_exit_it_1 ) : ( n184 ) ;
assign n186 =  ( n18 ) ? ( n182 ) : ( n185 ) ;
assign n187 =  ( n9 ) ? ( gb_exit_it_1 ) : ( n186 ) ;
assign n188 =  ( n4 ) ? ( gb_exit_it_1 ) : ( n187 ) ;
assign n189 =  ( n37 ) ? ( gb_exit_it_2 ) : ( gb_exit_it_2 ) ;
assign n190 =  ( n32 ) ? ( gb_exit_it_2 ) : ( n189 ) ;
assign n191 =  ( n25 ) ? ( gb_exit_it_2 ) : ( n190 ) ;
assign n192 =  ( n18 ) ? ( gb_exit_it_1 ) : ( n191 ) ;
assign n193 =  ( n9 ) ? ( gb_exit_it_2 ) : ( n192 ) ;
assign n194 =  ( n4 ) ? ( gb_exit_it_2 ) : ( n193 ) ;
assign n195 =  ( n37 ) ? ( gb_exit_it_3 ) : ( gb_exit_it_3 ) ;
assign n196 =  ( n32 ) ? ( gb_exit_it_3 ) : ( n195 ) ;
assign n197 =  ( n25 ) ? ( gb_exit_it_3 ) : ( n196 ) ;
assign n198 =  ( n18 ) ? ( gb_exit_it_2 ) : ( n197 ) ;
assign n199 =  ( n9 ) ? ( gb_exit_it_3 ) : ( n198 ) ;
assign n200 =  ( n4 ) ? ( gb_exit_it_3 ) : ( n199 ) ;
assign n201 =  ( n37 ) ? ( gb_exit_it_4 ) : ( gb_exit_it_4 ) ;
assign n202 =  ( n32 ) ? ( gb_exit_it_4 ) : ( n201 ) ;
assign n203 =  ( n25 ) ? ( gb_exit_it_4 ) : ( n202 ) ;
assign n204 =  ( n18 ) ? ( gb_exit_it_3 ) : ( n203 ) ;
assign n205 =  ( n9 ) ? ( gb_exit_it_4 ) : ( n204 ) ;
assign n206 =  ( n4 ) ? ( gb_exit_it_4 ) : ( n205 ) ;
assign n207 =  ( n37 ) ? ( gb_exit_it_5 ) : ( gb_exit_it_5 ) ;
assign n208 =  ( n32 ) ? ( gb_exit_it_5 ) : ( n207 ) ;
assign n209 =  ( n25 ) ? ( gb_exit_it_5 ) : ( n208 ) ;
assign n210 =  ( n18 ) ? ( gb_exit_it_4 ) : ( n209 ) ;
assign n211 =  ( n9 ) ? ( gb_exit_it_5 ) : ( n210 ) ;
assign n212 =  ( n4 ) ? ( gb_exit_it_5 ) : ( n211 ) ;
assign n213 =  ( n37 ) ? ( gb_exit_it_6 ) : ( gb_exit_it_6 ) ;
assign n214 =  ( n32 ) ? ( gb_exit_it_6 ) : ( n213 ) ;
assign n215 =  ( n25 ) ? ( gb_exit_it_6 ) : ( n214 ) ;
assign n216 =  ( n18 ) ? ( gb_exit_it_5 ) : ( n215 ) ;
assign n217 =  ( n9 ) ? ( gb_exit_it_6 ) : ( n216 ) ;
assign n218 =  ( n4 ) ? ( gb_exit_it_6 ) : ( n217 ) ;
assign n219 =  ( n37 ) ? ( gb_exit_it_7 ) : ( gb_exit_it_7 ) ;
assign n220 =  ( n32 ) ? ( gb_exit_it_7 ) : ( n219 ) ;
assign n221 =  ( n25 ) ? ( gb_exit_it_7 ) : ( n220 ) ;
assign n222 =  ( n18 ) ? ( gb_exit_it_6 ) : ( n221 ) ;
assign n223 =  ( n9 ) ? ( gb_exit_it_7 ) : ( n222 ) ;
assign n224 =  ( n4 ) ? ( gb_exit_it_7 ) : ( n223 ) ;
assign n225 =  ( n37 ) ? ( gb_exit_it_8 ) : ( gb_exit_it_8 ) ;
assign n226 =  ( n32 ) ? ( gb_exit_it_8 ) : ( n225 ) ;
assign n227 =  ( n25 ) ? ( gb_exit_it_8 ) : ( n226 ) ;
assign n228 =  ( n18 ) ? ( gb_exit_it_7 ) : ( n227 ) ;
assign n229 =  ( n9 ) ? ( gb_exit_it_8 ) : ( n228 ) ;
assign n230 =  ( n4 ) ? ( gb_exit_it_8 ) : ( n229 ) ;
assign n231 =  ( gb_p_cnt ) < ( 19'd307200 )  ;
assign n232 =  ( n231 ) ? ( n180 ) : ( 19'd307200 ) ;
assign n233 =  ( n37 ) ? ( gb_p_cnt ) : ( gb_p_cnt ) ;
assign n234 =  ( n32 ) ? ( gb_p_cnt ) : ( n233 ) ;
assign n235 =  ( n25 ) ? ( gb_p_cnt ) : ( n234 ) ;
assign n236 =  ( n18 ) ? ( n232 ) : ( n235 ) ;
assign n237 =  ( n9 ) ? ( gb_p_cnt ) : ( n236 ) ;
assign n238 =  ( n4 ) ? ( gb_p_cnt ) : ( n237 ) ;
assign n239 =  ( n37 ) ? ( gb_pp_it_1 ) : ( gb_pp_it_1 ) ;
assign n240 =  ( n32 ) ? ( gb_pp_it_1 ) : ( n239 ) ;
assign n241 =  ( n25 ) ? ( gb_pp_it_1 ) : ( n240 ) ;
assign n242 =  ( n18 ) ? ( 1'd1 ) : ( n241 ) ;
assign n243 =  ( n9 ) ? ( gb_pp_it_1 ) : ( n242 ) ;
assign n244 =  ( n4 ) ? ( gb_pp_it_1 ) : ( n243 ) ;
assign n245 =  ( n37 ) ? ( gb_pp_it_2 ) : ( gb_pp_it_2 ) ;
assign n246 =  ( n32 ) ? ( gb_pp_it_2 ) : ( n245 ) ;
assign n247 =  ( n25 ) ? ( gb_pp_it_2 ) : ( n246 ) ;
assign n248 =  ( n18 ) ? ( gb_pp_it_1 ) : ( n247 ) ;
assign n249 =  ( n9 ) ? ( gb_pp_it_2 ) : ( n248 ) ;
assign n250 =  ( n4 ) ? ( gb_pp_it_2 ) : ( n249 ) ;
assign n251 =  ( n37 ) ? ( gb_pp_it_3 ) : ( gb_pp_it_3 ) ;
assign n252 =  ( n32 ) ? ( gb_pp_it_3 ) : ( n251 ) ;
assign n253 =  ( n25 ) ? ( gb_pp_it_3 ) : ( n252 ) ;
assign n254 =  ( n18 ) ? ( gb_pp_it_2 ) : ( n253 ) ;
assign n255 =  ( n9 ) ? ( gb_pp_it_3 ) : ( n254 ) ;
assign n256 =  ( n4 ) ? ( gb_pp_it_3 ) : ( n255 ) ;
assign n257 =  ( n37 ) ? ( gb_pp_it_4 ) : ( gb_pp_it_4 ) ;
assign n258 =  ( n32 ) ? ( gb_pp_it_4 ) : ( n257 ) ;
assign n259 =  ( n25 ) ? ( gb_pp_it_4 ) : ( n258 ) ;
assign n260 =  ( n18 ) ? ( gb_pp_it_3 ) : ( n259 ) ;
assign n261 =  ( n9 ) ? ( gb_pp_it_4 ) : ( n260 ) ;
assign n262 =  ( n4 ) ? ( gb_pp_it_4 ) : ( n261 ) ;
assign n263 =  ( n37 ) ? ( gb_pp_it_5 ) : ( gb_pp_it_5 ) ;
assign n264 =  ( n32 ) ? ( gb_pp_it_5 ) : ( n263 ) ;
assign n265 =  ( n25 ) ? ( gb_pp_it_5 ) : ( n264 ) ;
assign n266 =  ( n18 ) ? ( gb_pp_it_4 ) : ( n265 ) ;
assign n267 =  ( n9 ) ? ( gb_pp_it_5 ) : ( n266 ) ;
assign n268 =  ( n4 ) ? ( gb_pp_it_5 ) : ( n267 ) ;
assign n269 =  ( n37 ) ? ( gb_pp_it_6 ) : ( gb_pp_it_6 ) ;
assign n270 =  ( n32 ) ? ( gb_pp_it_6 ) : ( n269 ) ;
assign n271 =  ( n25 ) ? ( gb_pp_it_6 ) : ( n270 ) ;
assign n272 =  ( n18 ) ? ( gb_pp_it_5 ) : ( n271 ) ;
assign n273 =  ( n9 ) ? ( gb_pp_it_6 ) : ( n272 ) ;
assign n274 =  ( n4 ) ? ( gb_pp_it_6 ) : ( n273 ) ;
assign n275 =  ( n37 ) ? ( gb_pp_it_7 ) : ( gb_pp_it_7 ) ;
assign n276 =  ( n32 ) ? ( gb_pp_it_7 ) : ( n275 ) ;
assign n277 =  ( n25 ) ? ( gb_pp_it_7 ) : ( n276 ) ;
assign n278 =  ( n18 ) ? ( gb_pp_it_6 ) : ( n277 ) ;
assign n279 =  ( n9 ) ? ( gb_pp_it_7 ) : ( n278 ) ;
assign n280 =  ( n4 ) ? ( gb_pp_it_7 ) : ( n279 ) ;
assign n281 =  ( n37 ) ? ( gb_pp_it_8 ) : ( gb_pp_it_8 ) ;
assign n282 =  ( n32 ) ? ( gb_pp_it_8 ) : ( n281 ) ;
assign n283 =  ( n25 ) ? ( gb_pp_it_8 ) : ( n282 ) ;
assign n284 =  ( n18 ) ? ( gb_pp_it_7 ) : ( n283 ) ;
assign n285 =  ( n9 ) ? ( gb_pp_it_8 ) : ( n284 ) ;
assign n286 =  ( n4 ) ? ( gb_pp_it_8 ) : ( n285 ) ;
assign n287 =  ( n37 ) ? ( gb_pp_it_9 ) : ( gb_pp_it_9 ) ;
assign n288 =  ( n32 ) ? ( gb_pp_it_9 ) : ( n287 ) ;
assign n289 =  ( n25 ) ? ( gb_pp_it_9 ) : ( n288 ) ;
assign n290 =  ( n18 ) ? ( gb_pp_it_8 ) : ( n289 ) ;
assign n291 =  ( n9 ) ? ( gb_pp_it_9 ) : ( n290 ) ;
assign n292 =  ( n4 ) ? ( gb_pp_it_9 ) : ( n291 ) ;
assign n293 =  ( n37 ) ? ( LB1D_buff ) : ( in_stream_buff_0 ) ;
assign n294 =  ( n32 ) ? ( in_stream_buff_0 ) : ( n293 ) ;
assign n295 =  ( n25 ) ? ( in_stream_buff_0 ) : ( n294 ) ;
assign n296 =  ( n18 ) ? ( in_stream_buff_0 ) : ( n295 ) ;
assign n297 =  ( n9 ) ? ( in_stream_buff_0 ) : ( n296 ) ;
assign n298 =  ( n4 ) ? ( in_stream_buff_0 ) : ( n297 ) ;
assign n299 =  ( n37 ) ? ( in_stream_buff_0 ) : ( in_stream_buff_1 ) ;
assign n300 =  ( n32 ) ? ( in_stream_buff_1 ) : ( n299 ) ;
assign n301 =  ( n25 ) ? ( in_stream_buff_1 ) : ( n300 ) ;
assign n302 =  ( n18 ) ? ( in_stream_buff_1 ) : ( n301 ) ;
assign n303 =  ( n9 ) ? ( in_stream_buff_1 ) : ( n302 ) ;
assign n304 =  ( n4 ) ? ( in_stream_buff_1 ) : ( n303 ) ;
assign n305 =  ( in_stream_full ) == ( 1'd1 )  ;
assign n306 =  ( n305 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n307 =  ( n37 ) ? ( 1'd0 ) : ( in_stream_empty ) ;
assign n308 =  ( n32 ) ? ( n306 ) : ( n307 ) ;
assign n309 =  ( n25 ) ? ( in_stream_empty ) : ( n308 ) ;
assign n310 =  ( n18 ) ? ( in_stream_empty ) : ( n309 ) ;
assign n311 =  ( n9 ) ? ( in_stream_empty ) : ( n310 ) ;
assign n312 =  ( n4 ) ? ( in_stream_empty ) : ( n311 ) ;
assign n313 =  ( in_stream_empty ) == ( 1'd1 )  ;
assign n314 =  ( n313 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n315 =  ( n37 ) ? ( n314 ) : ( in_stream_full ) ;
assign n316 =  ( n32 ) ? ( 1'd0 ) : ( n315 ) ;
assign n317 =  ( n25 ) ? ( in_stream_full ) : ( n316 ) ;
assign n318 =  ( n18 ) ? ( in_stream_full ) : ( n317 ) ;
assign n319 =  ( n9 ) ? ( in_stream_full ) : ( n318 ) ;
assign n320 =  ( n4 ) ? ( in_stream_full ) : ( n319 ) ;
assign n321 =  ( n305 ) ? ( in_stream_buff_1 ) : ( in_stream_buff_0 ) ;
assign n322 =  ( LB2D_proc_w ) == ( 64'd0 )  ;
assign n323 =  (  LB2D_proc_7 [ LB2D_proc_x ] )  ;
assign n324 =  ( LB2D_proc_w ) == ( 64'd1 )  ;
assign n325 =  (  LB2D_proc_0 [ LB2D_proc_x ] )  ;
assign n326 =  ( LB2D_proc_w ) == ( 64'd2 )  ;
assign n327 =  (  LB2D_proc_1 [ LB2D_proc_x ] )  ;
assign n328 =  ( LB2D_proc_w ) == ( 64'd3 )  ;
assign n329 =  (  LB2D_proc_2 [ LB2D_proc_x ] )  ;
assign n330 =  ( LB2D_proc_w ) == ( 64'd4 )  ;
assign n331 =  (  LB2D_proc_3 [ LB2D_proc_x ] )  ;
assign n332 =  ( LB2D_proc_w ) == ( 64'd5 )  ;
assign n333 =  (  LB2D_proc_4 [ LB2D_proc_x ] )  ;
assign n334 =  ( LB2D_proc_w ) == ( 64'd6 )  ;
assign n335 =  (  LB2D_proc_5 [ LB2D_proc_x ] )  ;
assign n336 =  (  LB2D_proc_6 [ LB2D_proc_x ] )  ;
assign n337 =  ( n334 ) ? ( n335 ) : ( n336 ) ;
assign n338 =  ( n332 ) ? ( n333 ) : ( n337 ) ;
assign n339 =  ( n330 ) ? ( n331 ) : ( n338 ) ;
assign n340 =  ( n328 ) ? ( n329 ) : ( n339 ) ;
assign n341 =  ( n326 ) ? ( n327 ) : ( n340 ) ;
assign n342 =  ( n324 ) ? ( n325 ) : ( n341 ) ;
assign n343 =  ( n322 ) ? ( n323 ) : ( n342 ) ;
assign n344 =  ( n334 ) ? ( n333 ) : ( n335 ) ;
assign n345 =  ( n332 ) ? ( n331 ) : ( n344 ) ;
assign n346 =  ( n330 ) ? ( n329 ) : ( n345 ) ;
assign n347 =  ( n328 ) ? ( n327 ) : ( n346 ) ;
assign n348 =  ( n326 ) ? ( n325 ) : ( n347 ) ;
assign n349 =  ( n324 ) ? ( n323 ) : ( n348 ) ;
assign n350 =  ( n322 ) ? ( n336 ) : ( n349 ) ;
assign n351 =  ( n334 ) ? ( n331 ) : ( n333 ) ;
assign n352 =  ( n332 ) ? ( n329 ) : ( n351 ) ;
assign n353 =  ( n330 ) ? ( n327 ) : ( n352 ) ;
assign n354 =  ( n328 ) ? ( n325 ) : ( n353 ) ;
assign n355 =  ( n326 ) ? ( n323 ) : ( n354 ) ;
assign n356 =  ( n324 ) ? ( n336 ) : ( n355 ) ;
assign n357 =  ( n322 ) ? ( n335 ) : ( n356 ) ;
assign n358 =  ( n334 ) ? ( n329 ) : ( n331 ) ;
assign n359 =  ( n332 ) ? ( n327 ) : ( n358 ) ;
assign n360 =  ( n330 ) ? ( n325 ) : ( n359 ) ;
assign n361 =  ( n328 ) ? ( n323 ) : ( n360 ) ;
assign n362 =  ( n326 ) ? ( n336 ) : ( n361 ) ;
assign n363 =  ( n324 ) ? ( n335 ) : ( n362 ) ;
assign n364 =  ( n322 ) ? ( n333 ) : ( n363 ) ;
assign n365 =  ( n334 ) ? ( n327 ) : ( n329 ) ;
assign n366 =  ( n332 ) ? ( n325 ) : ( n365 ) ;
assign n367 =  ( n330 ) ? ( n323 ) : ( n366 ) ;
assign n368 =  ( n328 ) ? ( n336 ) : ( n367 ) ;
assign n369 =  ( n326 ) ? ( n335 ) : ( n368 ) ;
assign n370 =  ( n324 ) ? ( n333 ) : ( n369 ) ;
assign n371 =  ( n322 ) ? ( n331 ) : ( n370 ) ;
assign n372 =  ( n334 ) ? ( n325 ) : ( n327 ) ;
assign n373 =  ( n332 ) ? ( n323 ) : ( n372 ) ;
assign n374 =  ( n330 ) ? ( n336 ) : ( n373 ) ;
assign n375 =  ( n328 ) ? ( n335 ) : ( n374 ) ;
assign n376 =  ( n326 ) ? ( n333 ) : ( n375 ) ;
assign n377 =  ( n324 ) ? ( n331 ) : ( n376 ) ;
assign n378 =  ( n322 ) ? ( n329 ) : ( n377 ) ;
assign n379 =  ( n334 ) ? ( n323 ) : ( n325 ) ;
assign n380 =  ( n332 ) ? ( n336 ) : ( n379 ) ;
assign n381 =  ( n330 ) ? ( n335 ) : ( n380 ) ;
assign n382 =  ( n328 ) ? ( n333 ) : ( n381 ) ;
assign n383 =  ( n326 ) ? ( n331 ) : ( n382 ) ;
assign n384 =  ( n324 ) ? ( n329 ) : ( n383 ) ;
assign n385 =  ( n322 ) ? ( n327 ) : ( n384 ) ;
assign n386 =  ( n334 ) ? ( n336 ) : ( n323 ) ;
assign n387 =  ( n332 ) ? ( n335 ) : ( n386 ) ;
assign n388 =  ( n330 ) ? ( n333 ) : ( n387 ) ;
assign n389 =  ( n328 ) ? ( n331 ) : ( n388 ) ;
assign n390 =  ( n326 ) ? ( n329 ) : ( n389 ) ;
assign n391 =  ( n324 ) ? ( n327 ) : ( n390 ) ;
assign n392 =  ( n322 ) ? ( n325 ) : ( n391 ) ;
assign n393 =  { ( n385 ) , ( n392 ) }  ;
assign n394 =  { ( n378 ) , ( n393 ) }  ;
assign n395 =  { ( n371 ) , ( n394 ) }  ;
assign n396 =  { ( n364 ) , ( n395 ) }  ;
assign n397 =  { ( n357 ) , ( n396 ) }  ;
assign n398 =  { ( n350 ) , ( n397 ) }  ;
assign n399 =  { ( n343 ) , ( n398 ) }  ;
assign n400 =  { ( n321 ) , ( n399 ) }  ;
assign n401 =  ( n30 ) ? ( slice_stream_buff_0 ) : ( n400 ) ;
assign n402 =  ( n37 ) ? ( slice_stream_buff_0 ) : ( slice_stream_buff_0 ) ;
assign n403 =  ( n32 ) ? ( n401 ) : ( n402 ) ;
assign n404 =  ( n25 ) ? ( slice_stream_buff_0 ) : ( n403 ) ;
assign n405 =  ( n18 ) ? ( slice_stream_buff_0 ) : ( n404 ) ;
assign n406 =  ( n9 ) ? ( slice_stream_buff_0 ) : ( n405 ) ;
assign n407 =  ( n4 ) ? ( slice_stream_buff_0 ) : ( n406 ) ;
assign n408 =  ( n30 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n409 =  ( n37 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_1 ) ;
assign n410 =  ( n32 ) ? ( n408 ) : ( n409 ) ;
assign n411 =  ( n25 ) ? ( slice_stream_buff_1 ) : ( n410 ) ;
assign n412 =  ( n18 ) ? ( slice_stream_buff_1 ) : ( n411 ) ;
assign n413 =  ( n9 ) ? ( slice_stream_buff_1 ) : ( n412 ) ;
assign n414 =  ( n4 ) ? ( slice_stream_buff_1 ) : ( n413 ) ;
assign n415 =  ( n88 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n416 =  ( n30 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n417 =  ( n37 ) ? ( slice_stream_empty ) : ( slice_stream_empty ) ;
assign n418 =  ( n32 ) ? ( n416 ) : ( n417 ) ;
assign n419 =  ( n25 ) ? ( n415 ) : ( n418 ) ;
assign n420 =  ( n18 ) ? ( slice_stream_empty ) : ( n419 ) ;
assign n421 =  ( n9 ) ? ( slice_stream_empty ) : ( n420 ) ;
assign n422 =  ( n4 ) ? ( slice_stream_empty ) : ( n421 ) ;
assign n423 =  ( slice_stream_empty ) == ( 1'd1 )  ;
assign n424 =  ( n423 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n425 =  ( n30 ) ? ( 1'd0 ) : ( n424 ) ;
assign n426 =  ( n37 ) ? ( slice_stream_full ) : ( slice_stream_full ) ;
assign n427 =  ( n32 ) ? ( n425 ) : ( n426 ) ;
assign n428 =  ( n25 ) ? ( 1'd0 ) : ( n427 ) ;
assign n429 =  ( n18 ) ? ( slice_stream_full ) : ( n428 ) ;
assign n430 =  ( n9 ) ? ( slice_stream_full ) : ( n429 ) ;
assign n431 =  ( n4 ) ? ( slice_stream_full ) : ( n430 ) ;
assign n432 =  ( LB2D_shift_x ) >= ( 9'd8 )  ;
assign n433 = n89[71:64] ;
assign n434 = LB2D_shift_0[71:64] ;
assign n435 = LB2D_shift_1[71:64] ;
assign n436 = LB2D_shift_2[71:64] ;
assign n437 = LB2D_shift_3[71:64] ;
assign n438 = LB2D_shift_4[71:64] ;
assign n439 = LB2D_shift_5[71:64] ;
assign n440 = LB2D_shift_6[71:64] ;
assign n441 = LB2D_shift_7[71:64] ;
assign n442 =  { ( n440 ) , ( n441 ) }  ;
assign n443 =  { ( n439 ) , ( n442 ) }  ;
assign n444 =  { ( n438 ) , ( n443 ) }  ;
assign n445 =  { ( n437 ) , ( n444 ) }  ;
assign n446 =  { ( n436 ) , ( n445 ) }  ;
assign n447 =  { ( n435 ) , ( n446 ) }  ;
assign n448 =  { ( n434 ) , ( n447 ) }  ;
assign n449 =  { ( n433 ) , ( n448 ) }  ;
assign n450 = n89[63:56] ;
assign n451 = LB2D_shift_0[63:56] ;
assign n452 = LB2D_shift_1[63:56] ;
assign n453 = LB2D_shift_2[63:56] ;
assign n454 = LB2D_shift_3[63:56] ;
assign n455 = LB2D_shift_4[63:56] ;
assign n456 = LB2D_shift_5[63:56] ;
assign n457 = LB2D_shift_6[63:56] ;
assign n458 = LB2D_shift_7[63:56] ;
assign n459 =  { ( n457 ) , ( n458 ) }  ;
assign n460 =  { ( n456 ) , ( n459 ) }  ;
assign n461 =  { ( n455 ) , ( n460 ) }  ;
assign n462 =  { ( n454 ) , ( n461 ) }  ;
assign n463 =  { ( n453 ) , ( n462 ) }  ;
assign n464 =  { ( n452 ) , ( n463 ) }  ;
assign n465 =  { ( n451 ) , ( n464 ) }  ;
assign n466 =  { ( n450 ) , ( n465 ) }  ;
assign n467 = n89[55:48] ;
assign n468 = LB2D_shift_0[55:48] ;
assign n469 = LB2D_shift_1[55:48] ;
assign n470 = LB2D_shift_2[55:48] ;
assign n471 = LB2D_shift_3[55:48] ;
assign n472 = LB2D_shift_4[55:48] ;
assign n473 = LB2D_shift_5[55:48] ;
assign n474 = LB2D_shift_6[55:48] ;
assign n475 = LB2D_shift_7[55:48] ;
assign n476 =  { ( n474 ) , ( n475 ) }  ;
assign n477 =  { ( n473 ) , ( n476 ) }  ;
assign n478 =  { ( n472 ) , ( n477 ) }  ;
assign n479 =  { ( n471 ) , ( n478 ) }  ;
assign n480 =  { ( n470 ) , ( n479 ) }  ;
assign n481 =  { ( n469 ) , ( n480 ) }  ;
assign n482 =  { ( n468 ) , ( n481 ) }  ;
assign n483 =  { ( n467 ) , ( n482 ) }  ;
assign n484 = n89[47:40] ;
assign n485 = LB2D_shift_0[47:40] ;
assign n486 = LB2D_shift_1[47:40] ;
assign n487 = LB2D_shift_2[47:40] ;
assign n488 = LB2D_shift_3[47:40] ;
assign n489 = LB2D_shift_4[47:40] ;
assign n490 = LB2D_shift_5[47:40] ;
assign n491 = LB2D_shift_6[47:40] ;
assign n492 = LB2D_shift_7[47:40] ;
assign n493 =  { ( n491 ) , ( n492 ) }  ;
assign n494 =  { ( n490 ) , ( n493 ) }  ;
assign n495 =  { ( n489 ) , ( n494 ) }  ;
assign n496 =  { ( n488 ) , ( n495 ) }  ;
assign n497 =  { ( n487 ) , ( n496 ) }  ;
assign n498 =  { ( n486 ) , ( n497 ) }  ;
assign n499 =  { ( n485 ) , ( n498 ) }  ;
assign n500 =  { ( n484 ) , ( n499 ) }  ;
assign n501 = n89[39:32] ;
assign n502 = LB2D_shift_0[39:32] ;
assign n503 = LB2D_shift_1[39:32] ;
assign n504 = LB2D_shift_2[39:32] ;
assign n505 = LB2D_shift_3[39:32] ;
assign n506 = LB2D_shift_4[39:32] ;
assign n507 = LB2D_shift_5[39:32] ;
assign n508 = LB2D_shift_6[39:32] ;
assign n509 = LB2D_shift_7[39:32] ;
assign n510 =  { ( n508 ) , ( n509 ) }  ;
assign n511 =  { ( n507 ) , ( n510 ) }  ;
assign n512 =  { ( n506 ) , ( n511 ) }  ;
assign n513 =  { ( n505 ) , ( n512 ) }  ;
assign n514 =  { ( n504 ) , ( n513 ) }  ;
assign n515 =  { ( n503 ) , ( n514 ) }  ;
assign n516 =  { ( n502 ) , ( n515 ) }  ;
assign n517 =  { ( n501 ) , ( n516 ) }  ;
assign n518 = n89[31:24] ;
assign n519 = LB2D_shift_0[31:24] ;
assign n520 = LB2D_shift_1[31:24] ;
assign n521 = LB2D_shift_2[31:24] ;
assign n522 = LB2D_shift_3[31:24] ;
assign n523 = LB2D_shift_4[31:24] ;
assign n524 = LB2D_shift_5[31:24] ;
assign n525 = LB2D_shift_6[31:24] ;
assign n526 = LB2D_shift_7[31:24] ;
assign n527 =  { ( n525 ) , ( n526 ) }  ;
assign n528 =  { ( n524 ) , ( n527 ) }  ;
assign n529 =  { ( n523 ) , ( n528 ) }  ;
assign n530 =  { ( n522 ) , ( n529 ) }  ;
assign n531 =  { ( n521 ) , ( n530 ) }  ;
assign n532 =  { ( n520 ) , ( n531 ) }  ;
assign n533 =  { ( n519 ) , ( n532 ) }  ;
assign n534 =  { ( n518 ) , ( n533 ) }  ;
assign n535 = n89[23:16] ;
assign n536 = LB2D_shift_0[23:16] ;
assign n537 = LB2D_shift_1[23:16] ;
assign n538 = LB2D_shift_2[23:16] ;
assign n539 = LB2D_shift_3[23:16] ;
assign n540 = LB2D_shift_4[23:16] ;
assign n541 = LB2D_shift_5[23:16] ;
assign n542 = LB2D_shift_6[23:16] ;
assign n543 = LB2D_shift_7[23:16] ;
assign n544 =  { ( n542 ) , ( n543 ) }  ;
assign n545 =  { ( n541 ) , ( n544 ) }  ;
assign n546 =  { ( n540 ) , ( n545 ) }  ;
assign n547 =  { ( n539 ) , ( n546 ) }  ;
assign n548 =  { ( n538 ) , ( n547 ) }  ;
assign n549 =  { ( n537 ) , ( n548 ) }  ;
assign n550 =  { ( n536 ) , ( n549 ) }  ;
assign n551 =  { ( n535 ) , ( n550 ) }  ;
assign n552 = n89[15:8] ;
assign n553 = LB2D_shift_0[15:8] ;
assign n554 = LB2D_shift_1[15:8] ;
assign n555 = LB2D_shift_2[15:8] ;
assign n556 = LB2D_shift_3[15:8] ;
assign n557 = LB2D_shift_4[15:8] ;
assign n558 = LB2D_shift_5[15:8] ;
assign n559 = LB2D_shift_6[15:8] ;
assign n560 = LB2D_shift_7[15:8] ;
assign n561 =  { ( n559 ) , ( n560 ) }  ;
assign n562 =  { ( n558 ) , ( n561 ) }  ;
assign n563 =  { ( n557 ) , ( n562 ) }  ;
assign n564 =  { ( n556 ) , ( n563 ) }  ;
assign n565 =  { ( n555 ) , ( n564 ) }  ;
assign n566 =  { ( n554 ) , ( n565 ) }  ;
assign n567 =  { ( n553 ) , ( n566 ) }  ;
assign n568 =  { ( n552 ) , ( n567 ) }  ;
assign n569 = n89[7:0] ;
assign n570 = LB2D_shift_0[7:0] ;
assign n571 = LB2D_shift_1[7:0] ;
assign n572 = LB2D_shift_2[7:0] ;
assign n573 = LB2D_shift_3[7:0] ;
assign n574 = LB2D_shift_4[7:0] ;
assign n575 = LB2D_shift_5[7:0] ;
assign n576 = LB2D_shift_6[7:0] ;
assign n577 = LB2D_shift_7[7:0] ;
assign n578 =  { ( n576 ) , ( n577 ) }  ;
assign n579 =  { ( n575 ) , ( n578 ) }  ;
assign n580 =  { ( n574 ) , ( n579 ) }  ;
assign n581 =  { ( n573 ) , ( n580 ) }  ;
assign n582 =  { ( n572 ) , ( n581 ) }  ;
assign n583 =  { ( n571 ) , ( n582 ) }  ;
assign n584 =  { ( n570 ) , ( n583 ) }  ;
assign n585 =  { ( n569 ) , ( n584 ) }  ;
assign n586 =  { ( n568 ) , ( n585 ) }  ;
assign n587 =  { ( n551 ) , ( n586 ) }  ;
assign n588 =  { ( n534 ) , ( n587 ) }  ;
assign n589 =  { ( n517 ) , ( n588 ) }  ;
assign n590 =  { ( n500 ) , ( n589 ) }  ;
assign n591 =  { ( n483 ) , ( n590 ) }  ;
assign n592 =  { ( n466 ) , ( n591 ) }  ;
assign n593 =  { ( n449 ) , ( n592 ) }  ;
assign n594 =  ( n432 ) ? ( n593 ) : ( stencil_stream_buff_0 ) ;
assign n595 =  ( n37 ) ? ( stencil_stream_buff_0 ) : ( stencil_stream_buff_0 ) ;
assign n596 =  ( n32 ) ? ( stencil_stream_buff_0 ) : ( n595 ) ;
assign n597 =  ( n25 ) ? ( n594 ) : ( n596 ) ;
assign n598 =  ( n18 ) ? ( stencil_stream_buff_0 ) : ( n597 ) ;
assign n599 =  ( n9 ) ? ( stencil_stream_buff_0 ) : ( n598 ) ;
assign n600 =  ( n4 ) ? ( stencil_stream_buff_0 ) : ( n599 ) ;
assign n601 =  ( n37 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_1 ) ;
assign n602 =  ( n32 ) ? ( stencil_stream_buff_1 ) : ( n601 ) ;
assign n603 =  ( n25 ) ? ( stencil_stream_buff_0 ) : ( n602 ) ;
assign n604 =  ( n18 ) ? ( stencil_stream_buff_1 ) : ( n603 ) ;
assign n605 =  ( n9 ) ? ( stencil_stream_buff_1 ) : ( n604 ) ;
assign n606 =  ( n4 ) ? ( stencil_stream_buff_1 ) : ( n605 ) ;
assign n607 =  ( n156 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n608 =  ( n23 ) ? ( stencil_stream_empty ) : ( 1'd0 ) ;
assign n609 =  ( n37 ) ? ( stencil_stream_empty ) : ( stencil_stream_empty ) ;
assign n610 =  ( n32 ) ? ( stencil_stream_empty ) : ( n609 ) ;
assign n611 =  ( n25 ) ? ( n608 ) : ( n610 ) ;
assign n612 =  ( n18 ) ? ( n607 ) : ( n611 ) ;
assign n613 =  ( n9 ) ? ( stencil_stream_empty ) : ( n612 ) ;
assign n614 =  ( n4 ) ? ( stencil_stream_empty ) : ( n613 ) ;
assign n615 =  ( n14 ) ? ( 1'd0 ) : ( 1'd0 ) ;
assign n616 =  ( stencil_stream_empty ) == ( 1'd1 )  ;
assign n617 =  ( n616 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n618 =  ( n23 ) ? ( stencil_stream_full ) : ( n617 ) ;
assign n619 =  ( n37 ) ? ( stencil_stream_full ) : ( stencil_stream_full ) ;
assign n620 =  ( n32 ) ? ( stencil_stream_full ) : ( n619 ) ;
assign n621 =  ( n25 ) ? ( n618 ) : ( n620 ) ;
assign n622 =  ( n18 ) ? ( n615 ) : ( n621 ) ;
assign n623 =  ( n9 ) ? ( stencil_stream_full ) : ( n622 ) ;
assign n624 =  ( n4 ) ? ( stencil_stream_full ) : ( n623 ) ;
assign n625 = ~ ( n4 ) ;
assign n626 = ~ ( n9 ) ;
assign n627 =  ( n625 ) & ( n626 )  ;
assign n628 = ~ ( n18 ) ;
assign n629 =  ( n627 ) & ( n628 )  ;
assign n630 = ~ ( n25 ) ;
assign n631 =  ( n629 ) & ( n630 )  ;
assign n632 = ~ ( n32 ) ;
assign n633 =  ( n631 ) & ( n632 )  ;
assign n634 = ~ ( n37 ) ;
assign n635 =  ( n633 ) & ( n634 )  ;
assign n636 =  ( n633 ) & ( n37 )  ;
assign n637 =  ( n631 ) & ( n32 )  ;
assign n638 = ~ ( n322 ) ;
assign n639 =  ( n637 ) & ( n638 )  ;
assign n640 =  ( n637 ) & ( n322 )  ;
assign n641 =  ( n629 ) & ( n25 )  ;
assign n642 =  ( n627 ) & ( n18 )  ;
assign n643 =  ( n625 ) & ( n9 )  ;
assign LB2D_proc_0_addr0 = n640 ? (LB2D_proc_x) : (0);
assign LB2D_proc_0_data0 = n640 ? (n321) : (LB2D_proc_0[0]);
assign n644 = ~ ( n324 ) ;
assign n645 =  ( n637 ) & ( n644 )  ;
assign n646 =  ( n637 ) & ( n324 )  ;
assign LB2D_proc_1_addr0 = n646 ? (LB2D_proc_x) : (0);
assign LB2D_proc_1_data0 = n646 ? (n321) : (LB2D_proc_1[0]);
assign n647 = ~ ( n326 ) ;
assign n648 =  ( n637 ) & ( n647 )  ;
assign n649 =  ( n637 ) & ( n326 )  ;
assign LB2D_proc_2_addr0 = n649 ? (LB2D_proc_x) : (0);
assign LB2D_proc_2_data0 = n649 ? (n321) : (LB2D_proc_2[0]);
assign n650 = ~ ( n328 ) ;
assign n651 =  ( n637 ) & ( n650 )  ;
assign n652 =  ( n637 ) & ( n328 )  ;
assign LB2D_proc_3_addr0 = n652 ? (LB2D_proc_x) : (0);
assign LB2D_proc_3_data0 = n652 ? (n321) : (LB2D_proc_3[0]);
assign n653 = ~ ( n330 ) ;
assign n654 =  ( n637 ) & ( n653 )  ;
assign n655 =  ( n637 ) & ( n330 )  ;
assign LB2D_proc_4_addr0 = n655 ? (LB2D_proc_x) : (0);
assign LB2D_proc_4_data0 = n655 ? (n321) : (LB2D_proc_4[0]);
assign n656 = ~ ( n332 ) ;
assign n657 =  ( n637 ) & ( n656 )  ;
assign n658 =  ( n637 ) & ( n332 )  ;
assign LB2D_proc_5_addr0 = n658 ? (LB2D_proc_x) : (0);
assign LB2D_proc_5_data0 = n658 ? (n321) : (LB2D_proc_5[0]);
assign n659 = ~ ( n334 ) ;
assign n660 =  ( n637 ) & ( n659 )  ;
assign n661 =  ( n637 ) & ( n334 )  ;
assign LB2D_proc_6_addr0 = n661 ? (LB2D_proc_x) : (0);
assign LB2D_proc_6_data0 = n661 ? (n321) : (LB2D_proc_6[0]);
assign n662 =  ( LB2D_proc_w ) == ( 64'd7 )  ;
assign n663 = ~ ( n662 ) ;
assign n664 =  ( n637 ) & ( n663 )  ;
assign n665 =  ( n637 ) & ( n662 )  ;
assign LB2D_proc_7_addr0 = n665 ? (LB2D_proc_x) : (0);
assign LB2D_proc_7_data0 = n665 ? (n321) : (LB2D_proc_7[0]);
/*
function [7:0] gb_fun ;
input [647:0] arg0;
    begin
//TODO: Add the specific function HERE.    end
endfunction
*/

always @(posedge clk) begin
   if(rst) begin
       LB1D_buff <= LB1D_buff;
       LB1D_it_1 <= LB1D_it_1;
       LB1D_p_cnt <= LB1D_p_cnt;
       LB2D_proc_w <= LB2D_proc_w;
       LB2D_proc_x <= LB2D_proc_x;
       LB2D_proc_y <= LB2D_proc_y;
       LB2D_shift_0 <= LB2D_shift_0;
       LB2D_shift_1 <= LB2D_shift_1;
       LB2D_shift_2 <= LB2D_shift_2;
       LB2D_shift_3 <= LB2D_shift_3;
       LB2D_shift_4 <= LB2D_shift_4;
       LB2D_shift_5 <= LB2D_shift_5;
       LB2D_shift_6 <= LB2D_shift_6;
       LB2D_shift_7 <= LB2D_shift_7;
       LB2D_shift_x <= LB2D_shift_x;
       LB2D_shift_y <= LB2D_shift_y;
       arg_0_TDATA <= arg_0_TDATA;
       arg_0_TVALID <= arg_0_TVALID;
       arg_1_TREADY <= arg_1_TREADY;
       gb_exit_it_1 <= gb_exit_it_1;
       gb_exit_it_2 <= gb_exit_it_2;
       gb_exit_it_3 <= gb_exit_it_3;
       gb_exit_it_4 <= gb_exit_it_4;
       gb_exit_it_5 <= gb_exit_it_5;
       gb_exit_it_6 <= gb_exit_it_6;
       gb_exit_it_7 <= gb_exit_it_7;
       gb_exit_it_8 <= gb_exit_it_8;
       gb_p_cnt <= gb_p_cnt;
       gb_pp_it_1 <= gb_pp_it_1;
       gb_pp_it_2 <= gb_pp_it_2;
       gb_pp_it_3 <= gb_pp_it_3;
       gb_pp_it_4 <= gb_pp_it_4;
       gb_pp_it_5 <= gb_pp_it_5;
       gb_pp_it_6 <= gb_pp_it_6;
       gb_pp_it_7 <= gb_pp_it_7;
       gb_pp_it_8 <= gb_pp_it_8;
       gb_pp_it_9 <= gb_pp_it_9;
       in_stream_buff_0 <= in_stream_buff_0;
       in_stream_buff_1 <= in_stream_buff_1;
       in_stream_empty <= in_stream_empty;
       in_stream_full <= in_stream_full;
       slice_stream_buff_0 <= slice_stream_buff_0;
       slice_stream_buff_1 <= slice_stream_buff_1;
       slice_stream_empty <= slice_stream_empty;
       slice_stream_full <= slice_stream_full;
       stencil_stream_buff_0 <= stencil_stream_buff_0;
       stencil_stream_buff_1 <= stencil_stream_buff_1;
       stencil_stream_empty <= stencil_stream_empty;
       stencil_stream_full <= stencil_stream_full;
   end
   else if(step) begin
       LB1D_buff <= n43;
       LB1D_it_1 <= n46;
       LB1D_p_cnt <= n57;
       LB2D_proc_w <= n68;
       LB2D_proc_x <= n79;
       LB2D_proc_y <= n87;
       LB2D_shift_0 <= n95;
       LB2D_shift_1 <= n101;
       LB2D_shift_2 <= n107;
       LB2D_shift_3 <= n113;
       LB2D_shift_4 <= n119;
       LB2D_shift_5 <= n125;
       LB2D_shift_6 <= n131;
       LB2D_shift_7 <= n137;
       LB2D_shift_x <= n144;
       LB2D_shift_y <= n155;
       arg_0_TDATA <= n164;
       arg_0_TVALID <= n172;
       arg_1_TREADY <= n179;
       gb_exit_it_1 <= n188;
       gb_exit_it_2 <= n194;
       gb_exit_it_3 <= n200;
       gb_exit_it_4 <= n206;
       gb_exit_it_5 <= n212;
       gb_exit_it_6 <= n218;
       gb_exit_it_7 <= n224;
       gb_exit_it_8 <= n230;
       gb_p_cnt <= n238;
       gb_pp_it_1 <= n244;
       gb_pp_it_2 <= n250;
       gb_pp_it_3 <= n256;
       gb_pp_it_4 <= n262;
       gb_pp_it_5 <= n268;
       gb_pp_it_6 <= n274;
       gb_pp_it_7 <= n280;
       gb_pp_it_8 <= n286;
       gb_pp_it_9 <= n292;
       in_stream_buff_0 <= n298;
       in_stream_buff_1 <= n304;
       in_stream_empty <= n312;
       in_stream_full <= n320;
       slice_stream_buff_0 <= n407;
       slice_stream_buff_1 <= n414;
       slice_stream_empty <= n422;
       slice_stream_full <= n431;
       stencil_stream_buff_0 <= n600;
       stencil_stream_buff_1 <= n606;
       stencil_stream_empty <= n614;
       stencil_stream_full <= n624;
       LB2D_proc_0 [ LB2D_proc_0_addr0 ] <= LB2D_proc_0_data0;
       LB2D_proc_1 [ LB2D_proc_1_addr0 ] <= LB2D_proc_1_data0;
       LB2D_proc_2 [ LB2D_proc_2_addr0 ] <= LB2D_proc_2_data0;
       LB2D_proc_3 [ LB2D_proc_3_addr0 ] <= LB2D_proc_3_data0;
       LB2D_proc_4 [ LB2D_proc_4_addr0 ] <= LB2D_proc_4_data0;
       LB2D_proc_5 [ LB2D_proc_5_addr0 ] <= LB2D_proc_5_data0;
       LB2D_proc_6 [ LB2D_proc_6_addr0 ] <= LB2D_proc_6_data0;
       LB2D_proc_7 [ LB2D_proc_7_addr0 ] <= LB2D_proc_7_data0;
   end
end
endmodule
