module SPEC_B(
arg_0_TREADY,
arg_1_TDATA,
arg_1_TVALID,
LB1D_buff,
LB1D_in,
LB1D_it_1,
LB1D_p_cnt,
LB1D_uIn,
LB2D_proc_w,
LB2D_proc_x,
LB2D_proc_y,
LB2D_shift_0,
LB2D_shift_1,
LB2D_shift_2,
LB2D_shift_3,
LB2D_shift_4,
LB2D_shift_5,
LB2D_shift_6,
LB2D_shift_7,
LB2D_shift_x,
LB2D_shift_y,
arg_0_TDATA,
arg_0_TVALID,
arg_1_TREADY,
gb_exit_it_1,
gb_exit_it_2,
gb_exit_it_3,
gb_exit_it_4,
gb_exit_it_5,
gb_exit_it_6,
gb_exit_it_7,
gb_exit_it_8,
gb_p_cnt,
gb_pp_it_1,
gb_pp_it_2,
gb_pp_it_3,
gb_pp_it_4,
gb_pp_it_5,
gb_pp_it_6,
gb_pp_it_7,
gb_pp_it_8,
gb_pp_it_9,
in_stream_buff_0,
in_stream_buff_1,
in_stream_empty,
in_stream_full,
slice_stream_buff_0,
slice_stream_buff_1,
slice_stream_empty,
slice_stream_full,
stencil_stream_buff_0,
stencil_stream_buff_1,
stencil_stream_empty,
stencil_stream_full,
clk,rst,
step
);
input            arg_0_TREADY;
input      [7:0] arg_1_TDATA;
input            arg_1_TVALID;
input clk;
input rst;
input step;
output      [7:0] LB1D_buff;
output      [7:0] LB1D_in;
output            LB1D_it_1;
output     [18:0] LB1D_p_cnt;
output      [7:0] LB1D_uIn;
output     [63:0] LB2D_proc_w;
output      [8:0] LB2D_proc_x;
output      [9:0] LB2D_proc_y;
output     [71:0] LB2D_shift_0;
output     [71:0] LB2D_shift_1;
output     [71:0] LB2D_shift_2;
output     [71:0] LB2D_shift_3;
output     [71:0] LB2D_shift_4;
output     [71:0] LB2D_shift_5;
output     [71:0] LB2D_shift_6;
output     [71:0] LB2D_shift_7;
output      [8:0] LB2D_shift_x;
output      [9:0] LB2D_shift_y;
output      [7:0] arg_0_TDATA;
output            arg_0_TVALID;
output            arg_1_TREADY;
output            gb_exit_it_1;
output            gb_exit_it_2;
output            gb_exit_it_3;
output            gb_exit_it_4;
output            gb_exit_it_5;
output            gb_exit_it_6;
output            gb_exit_it_7;
output            gb_exit_it_8;
output     [18:0] gb_p_cnt;
output            gb_pp_it_1;
output            gb_pp_it_2;
output            gb_pp_it_3;
output            gb_pp_it_4;
output            gb_pp_it_5;
output            gb_pp_it_6;
output            gb_pp_it_7;
output            gb_pp_it_8;
output            gb_pp_it_9;
output      [7:0] in_stream_buff_0;
output      [7:0] in_stream_buff_1;
output            in_stream_empty;
output            in_stream_full;
output     [71:0] slice_stream_buff_0;
output     [71:0] slice_stream_buff_1;
output            slice_stream_empty;
output            slice_stream_full;
output    [647:0] stencil_stream_buff_0;
output    [647:0] stencil_stream_buff_1;
output            stencil_stream_empty;
output            stencil_stream_full;
reg      [7:0] LB1D_buff;
reg      [7:0] LB1D_in;
reg            LB1D_it_1;
reg     [18:0] LB1D_p_cnt;
reg      [7:0] LB1D_uIn;
reg     [63:0] LB2D_proc_w;
reg      [8:0] LB2D_proc_x;
reg      [9:0] LB2D_proc_y;
reg     [71:0] LB2D_shift_0;
reg     [71:0] LB2D_shift_1;
reg     [71:0] LB2D_shift_2;
reg     [71:0] LB2D_shift_3;
reg     [71:0] LB2D_shift_4;
reg     [71:0] LB2D_shift_5;
reg     [71:0] LB2D_shift_6;
reg     [71:0] LB2D_shift_7;
reg      [8:0] LB2D_shift_x;
reg      [9:0] LB2D_shift_y;
reg      [7:0] arg_0_TDATA;
reg            arg_0_TVALID;
reg            arg_1_TREADY;
reg            gb_exit_it_1;
reg            gb_exit_it_2;
reg            gb_exit_it_3;
reg            gb_exit_it_4;
reg            gb_exit_it_5;
reg            gb_exit_it_6;
reg            gb_exit_it_7;
reg            gb_exit_it_8;
reg     [18:0] gb_p_cnt;
reg            gb_pp_it_1;
reg            gb_pp_it_2;
reg            gb_pp_it_3;
reg            gb_pp_it_4;
reg            gb_pp_it_5;
reg            gb_pp_it_6;
reg            gb_pp_it_7;
reg            gb_pp_it_8;
reg            gb_pp_it_9;
reg      [7:0] in_stream_buff_0;
reg      [7:0] in_stream_buff_1;
reg            in_stream_empty;
reg            in_stream_full;
reg     [71:0] slice_stream_buff_0;
reg     [71:0] slice_stream_buff_1;
reg            slice_stream_empty;
reg            slice_stream_full;
reg    [647:0] stencil_stream_buff_0;
reg    [647:0] stencil_stream_buff_1;
reg            stencil_stream_empty;
reg            stencil_stream_full;
wire            arg_0_TREADY;
wire      [7:0] arg_1_TDATA;
wire            arg_1_TVALID;
wire            n0;
wire            n1;
wire            n2;
wire            n3;
wire            n4;
wire            n5;
wire            n6;
wire            n7;
wire            n8;
wire            n9;
wire            n10;
wire            n11;
wire            n12;
wire            n13;
wire            n14;
wire            n15;
wire            n16;
wire            n17;
wire            n18;
wire            n19;
wire            n20;
wire            n21;
wire            n22;
wire            n23;
wire            n24;
wire            n25;
wire            n26;
wire            n27;
wire            n28;
wire            n29;
wire            n30;
wire            n31;
wire            n32;
wire            n33;
wire            n34;
wire            n35;
wire            n36;
wire            n37;
wire            n38;
wire      [7:0] n39;
wire      [7:0] n40;
wire      [7:0] n41;
wire      [7:0] n42;
wire      [7:0] n43;
wire      [7:0] n44;
wire      [7:0] n45;
wire      [7:0] n46;
wire      [7:0] n47;
wire      [7:0] n48;
wire      [7:0] n49;
wire      [7:0] n50;
wire      [7:0] n51;
wire      [7:0] n52;
wire     [18:0] n53;
wire            n54;
wire            n55;
wire            n56;
wire            n57;
wire            n58;
wire     [18:0] n59;
wire     [18:0] n60;
wire     [18:0] n61;
wire     [18:0] n62;
wire     [18:0] n63;
wire     [18:0] n64;
wire     [18:0] n65;
wire     [18:0] n66;
wire      [7:0] n67;
wire      [7:0] n68;
wire      [7:0] n69;
wire      [7:0] n70;
wire      [7:0] n71;
wire      [7:0] n72;
wire      [7:0] n73;
wire            n74;
wire            n75;
wire     [63:0] n76;
wire     [63:0] n77;
wire     [63:0] n78;
wire     [63:0] n79;
wire     [63:0] n80;
wire     [63:0] n81;
wire     [63:0] n82;
wire     [63:0] n83;
wire      [8:0] n84;
wire      [8:0] n85;
wire      [8:0] n86;
wire      [8:0] n87;
wire      [8:0] n88;
wire      [8:0] n89;
wire      [8:0] n90;
wire            n91;
wire      [9:0] n92;
wire      [9:0] n93;
wire      [9:0] n94;
wire      [9:0] n95;
wire      [9:0] n96;
wire      [9:0] n97;
wire      [9:0] n98;
wire      [9:0] n99;
wire     [71:0] n100;
wire     [71:0] n101;
wire     [71:0] n102;
wire     [71:0] n103;
wire     [71:0] n104;
wire     [71:0] n105;
wire     [71:0] n106;
wire     [71:0] n107;
wire     [71:0] n108;
wire     [71:0] n109;
wire     [71:0] n110;
wire     [71:0] n111;
wire     [71:0] n112;
wire     [71:0] n113;
wire     [71:0] n114;
wire     [71:0] n115;
wire     [71:0] n116;
wire     [71:0] n117;
wire     [71:0] n118;
wire     [71:0] n119;
wire     [71:0] n120;
wire     [71:0] n121;
wire     [71:0] n122;
wire     [71:0] n123;
wire     [71:0] n124;
wire     [71:0] n125;
wire     [71:0] n126;
wire     [71:0] n127;
wire     [71:0] n128;
wire     [71:0] n129;
wire     [71:0] n130;
wire     [71:0] n131;
wire     [71:0] n132;
wire     [71:0] n133;
wire     [71:0] n134;
wire            n135;
wire     [71:0] n136;
wire     [71:0] n137;
wire     [71:0] n138;
wire     [71:0] n139;
wire     [71:0] n140;
wire     [71:0] n141;
wire            n142;
wire            n143;
wire            n144;
wire            n145;
wire      [8:0] n146;
wire      [8:0] n147;
wire      [8:0] n148;
wire      [8:0] n149;
wire      [8:0] n150;
wire      [8:0] n151;
wire      [8:0] n152;
wire            n153;
wire            n154;
wire      [9:0] n155;
wire      [9:0] n156;
wire      [9:0] n157;
wire      [9:0] n158;
wire      [9:0] n159;
wire      [9:0] n160;
wire      [9:0] n161;
wire      [9:0] n162;
wire            n163;
wire    [647:0] n164;
wire      [7:0] n165;
wire      [7:0] n166;
wire      [7:0] n167;
wire      [7:0] n168;
wire      [7:0] n169;
wire      [7:0] n170;
wire      [7:0] n171;
wire            n172;
wire            n173;
wire            n174;
wire            n175;
wire            n176;
wire            n177;
wire            n178;
wire            n179;
wire            n180;
wire            n181;
wire            n182;
wire            n183;
wire            n184;
wire            n185;
wire            n186;
wire     [18:0] n187;
wire            n188;
wire            n189;
wire            n190;
wire            n191;
wire            n192;
wire            n193;
wire            n194;
wire            n195;
wire            n196;
wire            n197;
wire            n198;
wire            n199;
wire            n200;
wire            n201;
wire            n202;
wire            n203;
wire            n204;
wire            n205;
wire            n206;
wire            n207;
wire            n208;
wire            n209;
wire            n210;
wire            n211;
wire            n212;
wire            n213;
wire            n214;
wire            n215;
wire            n216;
wire            n217;
wire            n218;
wire            n219;
wire            n220;
wire            n221;
wire            n222;
wire            n223;
wire            n224;
wire            n225;
wire            n226;
wire            n227;
wire            n228;
wire            n229;
wire            n230;
wire     [18:0] n231;
wire     [18:0] n232;
wire     [18:0] n233;
wire     [18:0] n234;
wire     [18:0] n235;
wire     [18:0] n236;
wire            n237;
wire            n238;
wire            n239;
wire            n240;
wire            n241;
wire            n242;
wire            n243;
wire            n244;
wire            n245;
wire            n246;
wire            n247;
wire            n248;
wire            n249;
wire            n250;
wire            n251;
wire            n252;
wire            n253;
wire            n254;
wire            n255;
wire            n256;
wire            n257;
wire            n258;
wire            n259;
wire            n260;
wire            n261;
wire            n262;
wire            n263;
wire            n264;
wire            n265;
wire            n266;
wire            n267;
wire            n268;
wire            n269;
wire            n270;
wire            n271;
wire            n272;
wire            n273;
wire            n274;
wire            n275;
wire            n276;
wire            n277;
wire            n278;
wire            n279;
wire            n280;
wire            n281;
wire      [7:0] n282;
wire      [7:0] n283;
wire      [7:0] n284;
wire      [7:0] n285;
wire      [7:0] n286;
wire      [7:0] n287;
wire      [7:0] n288;
wire      [7:0] n289;
wire      [7:0] n290;
wire      [7:0] n291;
wire      [7:0] n292;
wire      [7:0] n293;
wire            n294;
wire            n295;
wire            n296;
wire            n297;
wire            n298;
wire            n299;
wire            n300;
wire            n301;
wire            n302;
wire            n303;
wire            n304;
wire            n305;
wire            n306;
wire            n307;
wire            n308;
wire            n309;
wire      [7:0] n310;
wire            n311;
wire      [8:0] n312;
wire      [7:0] n313;
wire            n314;
wire      [7:0] n315;
wire            n316;
wire      [7:0] n317;
wire            n318;
wire      [7:0] n319;
wire            n320;
wire      [7:0] n321;
wire            n322;
wire      [7:0] n323;
wire            n324;
wire      [7:0] n325;
wire      [7:0] n326;
wire      [7:0] n327;
wire      [7:0] n328;
wire      [7:0] n329;
wire      [7:0] n330;
wire      [7:0] n331;
wire      [7:0] n332;
wire      [7:0] n333;
wire      [7:0] n334;
wire      [7:0] n335;
wire      [7:0] n336;
wire      [7:0] n337;
wire      [7:0] n338;
wire      [7:0] n339;
wire      [7:0] n340;
wire      [7:0] n341;
wire      [7:0] n342;
wire      [7:0] n343;
wire      [7:0] n344;
wire      [7:0] n345;
wire      [7:0] n346;
wire      [7:0] n347;
wire      [7:0] n348;
wire      [7:0] n349;
wire      [7:0] n350;
wire      [7:0] n351;
wire      [7:0] n352;
wire      [7:0] n353;
wire      [7:0] n354;
wire      [7:0] n355;
wire      [7:0] n356;
wire      [7:0] n357;
wire      [7:0] n358;
wire      [7:0] n359;
wire      [7:0] n360;
wire      [7:0] n361;
wire      [7:0] n362;
wire      [7:0] n363;
wire      [7:0] n364;
wire      [7:0] n365;
wire      [7:0] n366;
wire      [7:0] n367;
wire      [7:0] n368;
wire      [7:0] n369;
wire      [7:0] n370;
wire      [7:0] n371;
wire      [7:0] n372;
wire      [7:0] n373;
wire      [7:0] n374;
wire      [7:0] n375;
wire      [7:0] n376;
wire      [7:0] n377;
wire      [7:0] n378;
wire      [7:0] n379;
wire      [7:0] n380;
wire      [7:0] n381;
wire      [7:0] n382;
wire     [15:0] n383;
wire     [23:0] n384;
wire     [31:0] n385;
wire     [39:0] n386;
wire     [47:0] n387;
wire     [55:0] n388;
wire     [63:0] n389;
wire     [71:0] n390;
wire     [71:0] n391;
wire     [71:0] n392;
wire     [71:0] n393;
wire     [71:0] n394;
wire     [71:0] n395;
wire     [71:0] n396;
wire     [71:0] n397;
wire     [71:0] n398;
wire     [71:0] n399;
wire     [71:0] n400;
wire     [71:0] n401;
wire     [71:0] n402;
wire            n403;
wire            n404;
wire            n405;
wire            n406;
wire            n407;
wire            n408;
wire            n409;
wire            n410;
wire            n411;
wire            n412;
wire            n413;
wire            n414;
wire            n415;
wire            n416;
wire            n417;
wire            n418;
wire            n419;
wire            n420;
wire      [7:0] n421;
wire      [7:0] n422;
wire      [7:0] n423;
wire      [7:0] n424;
wire      [7:0] n425;
wire      [7:0] n426;
wire      [7:0] n427;
wire      [7:0] n428;
wire      [7:0] n429;
wire     [15:0] n430;
wire     [23:0] n431;
wire     [31:0] n432;
wire     [39:0] n433;
wire     [47:0] n434;
wire     [55:0] n435;
wire     [63:0] n436;
wire     [71:0] n437;
wire      [7:0] n438;
wire      [7:0] n439;
wire      [7:0] n440;
wire      [7:0] n441;
wire      [7:0] n442;
wire      [7:0] n443;
wire      [7:0] n444;
wire      [7:0] n445;
wire      [7:0] n446;
wire     [15:0] n447;
wire     [23:0] n448;
wire     [31:0] n449;
wire     [39:0] n450;
wire     [47:0] n451;
wire     [55:0] n452;
wire     [63:0] n453;
wire     [71:0] n454;
wire      [7:0] n455;
wire      [7:0] n456;
wire      [7:0] n457;
wire      [7:0] n458;
wire      [7:0] n459;
wire      [7:0] n460;
wire      [7:0] n461;
wire      [7:0] n462;
wire      [7:0] n463;
wire     [15:0] n464;
wire     [23:0] n465;
wire     [31:0] n466;
wire     [39:0] n467;
wire     [47:0] n468;
wire     [55:0] n469;
wire     [63:0] n470;
wire     [71:0] n471;
wire      [7:0] n472;
wire      [7:0] n473;
wire      [7:0] n474;
wire      [7:0] n475;
wire      [7:0] n476;
wire      [7:0] n477;
wire      [7:0] n478;
wire      [7:0] n479;
wire      [7:0] n480;
wire     [15:0] n481;
wire     [23:0] n482;
wire     [31:0] n483;
wire     [39:0] n484;
wire     [47:0] n485;
wire     [55:0] n486;
wire     [63:0] n487;
wire     [71:0] n488;
wire      [7:0] n489;
wire      [7:0] n490;
wire      [7:0] n491;
wire      [7:0] n492;
wire      [7:0] n493;
wire      [7:0] n494;
wire      [7:0] n495;
wire      [7:0] n496;
wire      [7:0] n497;
wire     [15:0] n498;
wire     [23:0] n499;
wire     [31:0] n500;
wire     [39:0] n501;
wire     [47:0] n502;
wire     [55:0] n503;
wire     [63:0] n504;
wire     [71:0] n505;
wire      [7:0] n506;
wire      [7:0] n507;
wire      [7:0] n508;
wire      [7:0] n509;
wire      [7:0] n510;
wire      [7:0] n511;
wire      [7:0] n512;
wire      [7:0] n513;
wire      [7:0] n514;
wire     [15:0] n515;
wire     [23:0] n516;
wire     [31:0] n517;
wire     [39:0] n518;
wire     [47:0] n519;
wire     [55:0] n520;
wire     [63:0] n521;
wire     [71:0] n522;
wire      [7:0] n523;
wire      [7:0] n524;
wire      [7:0] n525;
wire      [7:0] n526;
wire      [7:0] n527;
wire      [7:0] n528;
wire      [7:0] n529;
wire      [7:0] n530;
wire      [7:0] n531;
wire     [15:0] n532;
wire     [23:0] n533;
wire     [31:0] n534;
wire     [39:0] n535;
wire     [47:0] n536;
wire     [55:0] n537;
wire     [63:0] n538;
wire     [71:0] n539;
wire      [7:0] n540;
wire      [7:0] n541;
wire      [7:0] n542;
wire      [7:0] n543;
wire      [7:0] n544;
wire      [7:0] n545;
wire      [7:0] n546;
wire      [7:0] n547;
wire      [7:0] n548;
wire     [15:0] n549;
wire     [23:0] n550;
wire     [31:0] n551;
wire     [39:0] n552;
wire     [47:0] n553;
wire     [55:0] n554;
wire     [63:0] n555;
wire     [71:0] n556;
wire      [7:0] n557;
wire      [7:0] n558;
wire      [7:0] n559;
wire      [7:0] n560;
wire      [7:0] n561;
wire      [7:0] n562;
wire      [7:0] n563;
wire      [7:0] n564;
wire      [7:0] n565;
wire     [15:0] n566;
wire     [23:0] n567;
wire     [31:0] n568;
wire     [39:0] n569;
wire     [47:0] n570;
wire     [55:0] n571;
wire     [63:0] n572;
wire     [71:0] n573;
wire    [143:0] n574;
wire    [215:0] n575;
wire    [287:0] n576;
wire    [359:0] n577;
wire    [431:0] n578;
wire    [503:0] n579;
wire    [575:0] n580;
wire    [647:0] n581;
wire    [647:0] n582;
wire    [647:0] n583;
wire    [647:0] n584;
wire    [647:0] n585;
wire    [647:0] n586;
wire    [647:0] n587;
wire    [647:0] n588;
wire    [647:0] n589;
wire    [647:0] n590;
wire    [647:0] n591;
wire    [647:0] n592;
wire            n593;
wire            n594;
wire            n595;
wire            n596;
wire            n597;
wire            n598;
wire            n599;
wire            n600;
wire            n601;
wire            n602;
wire            n603;
wire            n604;
wire            n605;
wire            n606;
wire            n607;
wire            n608;
wire            n609;
wire      [8:0] LB2D_proc_0_addr0;
wire      [7:0] LB2D_proc_0_data0;
wire            n610;
wire            n611;
wire            n612;
wire            n613;
wire            n614;
wire            n615;
wire            n616;
wire            n617;
wire            n618;
wire            n619;
wire            n620;
wire            n621;
wire            n622;
wire            n623;
wire            n624;
wire            n625;
wire      [8:0] LB2D_proc_1_addr0;
wire      [7:0] LB2D_proc_1_data0;
wire            n626;
wire            n627;
wire            n628;
wire      [8:0] LB2D_proc_2_addr0;
wire      [7:0] LB2D_proc_2_data0;
wire            n629;
wire            n630;
wire            n631;
wire      [8:0] LB2D_proc_3_addr0;
wire      [7:0] LB2D_proc_3_data0;
wire            n632;
wire            n633;
wire            n634;
wire      [8:0] LB2D_proc_4_addr0;
wire      [7:0] LB2D_proc_4_data0;
wire            n635;
wire            n636;
wire            n637;
wire      [8:0] LB2D_proc_5_addr0;
wire      [7:0] LB2D_proc_5_data0;
wire            n638;
wire            n639;
wire            n640;
wire      [8:0] LB2D_proc_6_addr0;
wire      [7:0] LB2D_proc_6_data0;
wire            n641;
wire            n642;
wire            n643;
wire      [8:0] LB2D_proc_7_addr0;
wire      [7:0] LB2D_proc_7_data0;
wire            n644;
wire            n645;
wire            n646;
reg      [7:0] LB2D_proc_0[487:0];
reg      [7:0] LB2D_proc_1[487:0];
reg      [7:0] LB2D_proc_2[487:0];
reg      [7:0] LB2D_proc_3[487:0];
reg      [7:0] LB2D_proc_4[487:0];
reg      [7:0] LB2D_proc_5[487:0];
reg      [7:0] LB2D_proc_6[487:0];
reg      [7:0] LB2D_proc_7[487:0];
wire clk;
wire rst;
wire step;
assign n0 =  ( arg_1_TREADY ) == ( 1'd1 )  ;
assign n1 =  ( arg_1_TVALID ) == ( 1'd1 )  ;
assign n2 =  ( n0 ) & ( n1 )  ;
assign n3 =  ( arg_0_TREADY ) == ( 1'd0 )  ;
assign n4 =  ( n2 ) & ( n3 )  ;
assign n5 =  ( arg_0_TVALID ) == ( 1'd0 )  ;
assign n6 =  ( gb_exit_it_1 ) == ( 1'd0 )  ;
assign n7 =  ( stencil_stream_empty ) == ( 1'd0 )  ;
assign n8 =  ( n6 ) & ( n7 )  ;
assign n9 =  ( gb_exit_it_1 ) == ( 1'd1 )  ;
assign n10 =  ( gb_exit_it_8 ) == ( 1'd0 )  ;
assign n11 =  ( n9 ) & ( n10 )  ;
assign n12 =  ( n8 ) | ( n11 )  ;
assign n13 =  ( n5 ) & ( n12 )  ;
assign n14 =  ( slice_stream_empty ) == ( 1'd0 )  ;
assign n15 =  ( LB2D_shift_x ) != ( 9'd488 )  ;
assign n16 =  ( n14 ) & ( n15 )  ;
assign n17 =  ( stencil_stream_full ) == ( 1'd0 )  ;
assign n18 =  ( LB2D_shift_x ) < ( 9'd8 )  ;
assign n19 =  ( LB2D_shift_x ) > ( 9'd0 )  ;
assign n20 =  ( n18 ) & ( n19 )  ;
assign n21 =  ( n17 ) | ( n20 )  ;
assign n22 =  ( n16 ) & ( n21 )  ;
assign n23 =  ( in_stream_empty ) == ( 1'd0 )  ;
assign n24 =  ( slice_stream_full ) == ( 1'd0 )  ;
assign n25 =  ( LB2D_proc_y ) < ( 10'd8 )  ;
assign n26 =  ( n24 ) | ( n25 )  ;
assign n27 =  ( n23 ) & ( n26 )  ;
assign n28 =  ( in_stream_full ) == ( 1'd0 )  ;
assign n29 =  ( n0 ) & ( n28 )  ;
assign n30 =  ( LB1D_it_1 ) == ( 1'd0 )  ;
assign n31 =  ( n29 ) & ( n30 )  ;
assign n32 =  ( LB1D_p_cnt ) == ( 19'd316224 )  ;
assign n33 =  ( n31 ) & ( n32 )  ;
assign n34 =  ( arg_1_TREADY ) == ( 1'd0 )  ;
assign n35 =  ( n34 ) & ( n28 )  ;
assign n36 =  ( n35 ) & ( n30 )  ;
assign n37 =  ( LB1D_it_1 ) == ( 1'd1 )  ;
assign n38 =  ( n35 ) & ( n37 )  ;
assign n39 =  ( n38 ) ? ( LB1D_uIn ) : ( LB1D_buff ) ;
assign n40 =  ( n36 ) ? ( LB1D_uIn ) : ( n39 ) ;
assign n41 =  ( n33 ) ? ( LB1D_uIn ) : ( n40 ) ;
assign n42 =  ( n27 ) ? ( LB1D_buff ) : ( n41 ) ;
assign n43 =  ( n22 ) ? ( LB1D_buff ) : ( n42 ) ;
assign n44 =  ( n13 ) ? ( LB1D_buff ) : ( n43 ) ;
assign n45 =  ( n4 ) ? ( LB1D_buff ) : ( n44 ) ;
assign n46 =  ( n38 ) ? ( LB1D_in ) : ( LB1D_in ) ;
assign n47 =  ( n36 ) ? ( LB1D_in ) : ( n46 ) ;
assign n48 =  ( n33 ) ? ( LB1D_in ) : ( n47 ) ;
assign n49 =  ( n27 ) ? ( LB1D_in ) : ( n48 ) ;
assign n50 =  ( n22 ) ? ( LB1D_in ) : ( n49 ) ;
assign n51 =  ( n13 ) ? ( LB1D_in ) : ( n50 ) ;
assign n52 =  ( n4 ) ? ( arg_1_TDATA ) : ( n51 ) ;
assign n53 =  ( 19'd316224 ) - ( 19'd1 )  ;
assign n54 =  ( LB1D_p_cnt ) == ( n53 )  ;
assign n55 =  ( n54 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n56 =  ( n38 ) ? ( n55 ) : ( LB1D_it_1 ) ;
assign n57 =  ( n36 ) ? ( 1'd1 ) : ( n56 ) ;
assign n58 =  ( n33 ) ? ( 1'd0 ) : ( n57 ) ;
assign n59 =  ( LB1D_p_cnt ) + ( 19'd1 )  ;
assign n60 =  ( n38 ) ? ( n59 ) : ( LB1D_p_cnt ) ;
assign n61 =  ( n36 ) ? ( n59 ) : ( n60 ) ;
assign n62 =  ( n33 ) ? ( 19'd0 ) : ( n61 ) ;
assign n63 =  ( n27 ) ? ( LB1D_p_cnt ) : ( n62 ) ;
assign n64 =  ( n22 ) ? ( LB1D_p_cnt ) : ( n63 ) ;
assign n65 =  ( n13 ) ? ( LB1D_p_cnt ) : ( n64 ) ;
assign n66 =  ( n4 ) ? ( LB1D_p_cnt ) : ( n65 ) ;
assign n67 =  ( n38 ) ? ( LB1D_in ) : ( LB1D_uIn ) ;
assign n68 =  ( n36 ) ? ( LB1D_in ) : ( n67 ) ;
assign n69 =  ( n33 ) ? ( LB1D_in ) : ( n68 ) ;
assign n70 =  ( n27 ) ? ( LB1D_uIn ) : ( n69 ) ;
assign n71 =  ( n22 ) ? ( LB1D_uIn ) : ( n70 ) ;
assign n72 =  ( n13 ) ? ( LB1D_uIn ) : ( n71 ) ;
assign n73 =  ( n4 ) ? ( LB1D_uIn ) : ( n72 ) ;
assign n74 =  ( LB2D_proc_x ) == ( 9'd488 )  ;
assign n75 =  ( LB2D_proc_w ) == ( 64'd7 )  ;
assign n76 =  ( LB2D_proc_w ) + ( 64'd1 )  ;
assign n77 =  ( n75 ) ? ( 64'd0 ) : ( n76 ) ;
assign n78 =  ( n74 ) ? ( n77 ) : ( LB2D_proc_w ) ;
assign n79 =  ( n38 ) ? ( LB2D_proc_w ) : ( LB2D_proc_w ) ;
assign n80 =  ( n27 ) ? ( n78 ) : ( n79 ) ;
assign n81 =  ( n22 ) ? ( LB2D_proc_w ) : ( n80 ) ;
assign n82 =  ( n13 ) ? ( LB2D_proc_w ) : ( n81 ) ;
assign n83 =  ( n4 ) ? ( LB2D_proc_w ) : ( n82 ) ;
assign n84 =  ( LB2D_proc_x ) + ( 9'd1 )  ;
assign n85 =  ( n74 ) ? ( 9'd1 ) : ( n84 ) ;
assign n86 =  ( n38 ) ? ( LB2D_proc_x ) : ( LB2D_proc_x ) ;
assign n87 =  ( n27 ) ? ( n85 ) : ( n86 ) ;
assign n88 =  ( n22 ) ? ( LB2D_proc_x ) : ( n87 ) ;
assign n89 =  ( n13 ) ? ( LB2D_proc_x ) : ( n88 ) ;
assign n90 =  ( n4 ) ? ( LB2D_proc_x ) : ( n89 ) ;
assign n91 =  ( LB2D_proc_y ) == ( 10'd648 )  ;
assign n92 =  ( LB2D_proc_y ) + ( 10'd1 )  ;
assign n93 =  ( n91 ) ? ( 10'd0 ) : ( n92 ) ;
assign n94 =  ( n74 ) ? ( n93 ) : ( LB2D_proc_y ) ;
assign n95 =  ( n38 ) ? ( LB2D_proc_y ) : ( LB2D_proc_y ) ;
assign n96 =  ( n27 ) ? ( n94 ) : ( n95 ) ;
assign n97 =  ( n22 ) ? ( LB2D_proc_y ) : ( n96 ) ;
assign n98 =  ( n13 ) ? ( LB2D_proc_y ) : ( n97 ) ;
assign n99 =  ( n4 ) ? ( LB2D_proc_y ) : ( n98 ) ;
assign n100 =  ( n38 ) ? ( LB2D_shift_0 ) : ( LB2D_shift_0 ) ;
assign n101 =  ( n27 ) ? ( LB2D_shift_0 ) : ( n100 ) ;
assign n102 =  ( n22 ) ? ( LB2D_shift_1 ) : ( n101 ) ;
assign n103 =  ( n13 ) ? ( LB2D_shift_0 ) : ( n102 ) ;
assign n104 =  ( n4 ) ? ( LB2D_shift_0 ) : ( n103 ) ;
assign n105 =  ( n38 ) ? ( LB2D_shift_1 ) : ( LB2D_shift_1 ) ;
assign n106 =  ( n27 ) ? ( LB2D_shift_1 ) : ( n105 ) ;
assign n107 =  ( n22 ) ? ( LB2D_shift_2 ) : ( n106 ) ;
assign n108 =  ( n13 ) ? ( LB2D_shift_1 ) : ( n107 ) ;
assign n109 =  ( n4 ) ? ( LB2D_shift_1 ) : ( n108 ) ;
assign n110 =  ( n38 ) ? ( LB2D_shift_2 ) : ( LB2D_shift_2 ) ;
assign n111 =  ( n27 ) ? ( LB2D_shift_2 ) : ( n110 ) ;
assign n112 =  ( n22 ) ? ( LB2D_shift_3 ) : ( n111 ) ;
assign n113 =  ( n13 ) ? ( LB2D_shift_2 ) : ( n112 ) ;
assign n114 =  ( n4 ) ? ( LB2D_shift_2 ) : ( n113 ) ;
assign n115 =  ( n38 ) ? ( LB2D_shift_3 ) : ( LB2D_shift_3 ) ;
assign n116 =  ( n27 ) ? ( LB2D_shift_3 ) : ( n115 ) ;
assign n117 =  ( n22 ) ? ( LB2D_shift_4 ) : ( n116 ) ;
assign n118 =  ( n13 ) ? ( LB2D_shift_3 ) : ( n117 ) ;
assign n119 =  ( n4 ) ? ( LB2D_shift_3 ) : ( n118 ) ;
assign n120 =  ( n38 ) ? ( LB2D_shift_4 ) : ( LB2D_shift_4 ) ;
assign n121 =  ( n27 ) ? ( LB2D_shift_4 ) : ( n120 ) ;
assign n122 =  ( n22 ) ? ( LB2D_shift_5 ) : ( n121 ) ;
assign n123 =  ( n13 ) ? ( LB2D_shift_4 ) : ( n122 ) ;
assign n124 =  ( n4 ) ? ( LB2D_shift_4 ) : ( n123 ) ;
assign n125 =  ( n38 ) ? ( LB2D_shift_5 ) : ( LB2D_shift_5 ) ;
assign n126 =  ( n27 ) ? ( LB2D_shift_5 ) : ( n125 ) ;
assign n127 =  ( n22 ) ? ( LB2D_shift_6 ) : ( n126 ) ;
assign n128 =  ( n13 ) ? ( LB2D_shift_5 ) : ( n127 ) ;
assign n129 =  ( n4 ) ? ( LB2D_shift_5 ) : ( n128 ) ;
assign n130 =  ( n38 ) ? ( LB2D_shift_6 ) : ( LB2D_shift_6 ) ;
assign n131 =  ( n27 ) ? ( LB2D_shift_6 ) : ( n130 ) ;
assign n132 =  ( n22 ) ? ( LB2D_shift_7 ) : ( n131 ) ;
assign n133 =  ( n13 ) ? ( LB2D_shift_6 ) : ( n132 ) ;
assign n134 =  ( n4 ) ? ( LB2D_shift_6 ) : ( n133 ) ;
assign n135 =  ( slice_stream_full ) == ( 1'd1 )  ;
assign n136 =  ( n135 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n137 =  ( n38 ) ? ( LB2D_shift_7 ) : ( LB2D_shift_7 ) ;
assign n138 =  ( n27 ) ? ( LB2D_shift_7 ) : ( n137 ) ;
assign n139 =  ( n22 ) ? ( n136 ) : ( n138 ) ;
assign n140 =  ( n13 ) ? ( LB2D_shift_7 ) : ( n139 ) ;
assign n141 =  ( n4 ) ? ( LB2D_shift_7 ) : ( n140 ) ;
assign n142 =  ( LB2D_shift_x ) == ( 9'd488 )  ;
assign n143 =  ( n14 ) & ( n142 )  ;
assign n144 =  ( n17 ) | ( n18 )  ;
assign n145 =  ( n143 ) & ( n144 )  ;
assign n146 =  ( LB2D_shift_x ) + ( 9'd1 )  ;
assign n147 =  ( n38 ) ? ( LB2D_shift_x ) : ( LB2D_shift_x ) ;
assign n148 =  ( n27 ) ? ( LB2D_shift_x ) : ( n147 ) ;
assign n149 =  ( n22 ) ? ( n146 ) : ( n148 ) ;
assign n150 =  ( n145 ) ? ( 9'd0 ) : ( n149 ) ;
assign n151 =  ( n13 ) ? ( LB2D_shift_x ) : ( n150 ) ;
assign n152 =  ( n4 ) ? ( LB2D_shift_x ) : ( n151 ) ;
assign n153 =  ( LB2D_shift_y ) < ( 10'd640 )  ;
assign n154 =  ( LB2D_shift_x ) < ( 9'd488 )  ;
assign n155 =  ( LB2D_shift_y ) + ( 10'd1 )  ;
assign n156 =  ( n154 ) ? ( LB2D_shift_y ) : ( n155 ) ;
assign n157 =  ( n153 ) ? ( n156 ) : ( 10'd640 ) ;
assign n158 =  ( n38 ) ? ( LB2D_shift_y ) : ( LB2D_shift_y ) ;
assign n159 =  ( n27 ) ? ( LB2D_shift_y ) : ( n158 ) ;
assign n160 =  ( n22 ) ? ( n157 ) : ( n159 ) ;
assign n161 =  ( n13 ) ? ( LB2D_shift_y ) : ( n160 ) ;
assign n162 =  ( n4 ) ? ( LB2D_shift_y ) : ( n161 ) ;
assign n163 =  ( stencil_stream_full ) == ( 1'd1 )  ;
assign n164 =  ( n163 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_0 ) ;
//assign n165 = gb_fun(n164) ;
gb_fun gb_fun_U (
        .a (n164),
        .b (n165)
        );

assign n166 =  ( n38 ) ? ( arg_0_TDATA ) : ( arg_0_TDATA ) ;
assign n167 =  ( n33 ) ? ( arg_0_TDATA ) : ( n166 ) ;
assign n168 =  ( n27 ) ? ( arg_0_TDATA ) : ( n167 ) ;
assign n169 =  ( n22 ) ? ( arg_0_TDATA ) : ( n168 ) ;
assign n170 =  ( n13 ) ? ( n165 ) : ( n169 ) ;
assign n171 =  ( n4 ) ? ( arg_0_TDATA ) : ( n170 ) ;
assign n172 =  ( gb_pp_it_8 ) == ( 1'd1 )  ;
assign n173 =  ( n172 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n174 =  ( n38 ) ? ( arg_0_TVALID ) : ( arg_0_TVALID ) ;
assign n175 =  ( n33 ) ? ( arg_0_TVALID ) : ( n174 ) ;
assign n176 =  ( n27 ) ? ( arg_0_TVALID ) : ( n175 ) ;
assign n177 =  ( n22 ) ? ( arg_0_TVALID ) : ( n176 ) ;
assign n178 =  ( n13 ) ? ( n173 ) : ( n177 ) ;
assign n179 =  ( n4 ) ? ( arg_0_TVALID ) : ( n178 ) ;
assign n180 =  ( n38 ) ? ( 1'd1 ) : ( arg_1_TREADY ) ;
assign n181 =  ( n36 ) ? ( 1'd1 ) : ( n180 ) ;
assign n182 =  ( n33 ) ? ( 1'd1 ) : ( n181 ) ;
assign n183 =  ( n27 ) ? ( arg_1_TREADY ) : ( n182 ) ;
assign n184 =  ( n22 ) ? ( arg_1_TREADY ) : ( n183 ) ;
assign n185 =  ( n13 ) ? ( arg_1_TREADY ) : ( n184 ) ;
assign n186 =  ( n4 ) ? ( 1'd0 ) : ( n185 ) ;
assign n187 =  ( gb_p_cnt ) + ( 19'd1 )  ;
assign n188 =  ( n187 ) == ( 19'd307200 )  ;
assign n189 =  ( n188 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n190 =  ( n38 ) ? ( gb_exit_it_1 ) : ( gb_exit_it_1 ) ;
assign n191 =  ( n27 ) ? ( gb_exit_it_1 ) : ( n190 ) ;
assign n192 =  ( n22 ) ? ( gb_exit_it_1 ) : ( n191 ) ;
assign n193 =  ( n13 ) ? ( n189 ) : ( n192 ) ;
assign n194 =  ( n4 ) ? ( gb_exit_it_1 ) : ( n193 ) ;
assign n195 =  ( n38 ) ? ( gb_exit_it_2 ) : ( gb_exit_it_2 ) ;
assign n196 =  ( n27 ) ? ( gb_exit_it_2 ) : ( n195 ) ;
assign n197 =  ( n22 ) ? ( gb_exit_it_2 ) : ( n196 ) ;
assign n198 =  ( n13 ) ? ( gb_exit_it_1 ) : ( n197 ) ;
assign n199 =  ( n4 ) ? ( gb_exit_it_2 ) : ( n198 ) ;
assign n200 =  ( n38 ) ? ( gb_exit_it_3 ) : ( gb_exit_it_3 ) ;
assign n201 =  ( n27 ) ? ( gb_exit_it_3 ) : ( n200 ) ;
assign n202 =  ( n22 ) ? ( gb_exit_it_3 ) : ( n201 ) ;
assign n203 =  ( n13 ) ? ( gb_exit_it_2 ) : ( n202 ) ;
assign n204 =  ( n4 ) ? ( gb_exit_it_3 ) : ( n203 ) ;
assign n205 =  ( n38 ) ? ( gb_exit_it_4 ) : ( gb_exit_it_4 ) ;
assign n206 =  ( n27 ) ? ( gb_exit_it_4 ) : ( n205 ) ;
assign n207 =  ( n22 ) ? ( gb_exit_it_4 ) : ( n206 ) ;
assign n208 =  ( n13 ) ? ( gb_exit_it_3 ) : ( n207 ) ;
assign n209 =  ( n4 ) ? ( gb_exit_it_4 ) : ( n208 ) ;
assign n210 =  ( n38 ) ? ( gb_exit_it_5 ) : ( gb_exit_it_5 ) ;
assign n211 =  ( n27 ) ? ( gb_exit_it_5 ) : ( n210 ) ;
assign n212 =  ( n22 ) ? ( gb_exit_it_5 ) : ( n211 ) ;
assign n213 =  ( n13 ) ? ( gb_exit_it_4 ) : ( n212 ) ;
assign n214 =  ( n4 ) ? ( gb_exit_it_5 ) : ( n213 ) ;
assign n215 =  ( n38 ) ? ( gb_exit_it_6 ) : ( gb_exit_it_6 ) ;
assign n216 =  ( n27 ) ? ( gb_exit_it_6 ) : ( n215 ) ;
assign n217 =  ( n22 ) ? ( gb_exit_it_6 ) : ( n216 ) ;
assign n218 =  ( n13 ) ? ( gb_exit_it_5 ) : ( n217 ) ;
assign n219 =  ( n4 ) ? ( gb_exit_it_6 ) : ( n218 ) ;
assign n220 =  ( n38 ) ? ( gb_exit_it_7 ) : ( gb_exit_it_7 ) ;
assign n221 =  ( n27 ) ? ( gb_exit_it_7 ) : ( n220 ) ;
assign n222 =  ( n22 ) ? ( gb_exit_it_7 ) : ( n221 ) ;
assign n223 =  ( n13 ) ? ( gb_exit_it_6 ) : ( n222 ) ;
assign n224 =  ( n4 ) ? ( gb_exit_it_7 ) : ( n223 ) ;
assign n225 =  ( n38 ) ? ( gb_exit_it_8 ) : ( gb_exit_it_8 ) ;
assign n226 =  ( n27 ) ? ( gb_exit_it_8 ) : ( n225 ) ;
assign n227 =  ( n22 ) ? ( gb_exit_it_8 ) : ( n226 ) ;
assign n228 =  ( n13 ) ? ( gb_exit_it_7 ) : ( n227 ) ;
assign n229 =  ( n4 ) ? ( gb_exit_it_8 ) : ( n228 ) ;
assign n230 =  ( gb_p_cnt ) < ( 19'd307200 )  ;
assign n231 =  ( n230 ) ? ( n187 ) : ( 19'd307200 ) ;
assign n232 =  ( n38 ) ? ( gb_p_cnt ) : ( gb_p_cnt ) ;
assign n233 =  ( n27 ) ? ( gb_p_cnt ) : ( n232 ) ;
assign n234 =  ( n22 ) ? ( gb_p_cnt ) : ( n233 ) ;
assign n235 =  ( n13 ) ? ( n231 ) : ( n234 ) ;
assign n236 =  ( n4 ) ? ( gb_p_cnt ) : ( n235 ) ;
assign n237 =  ( n38 ) ? ( gb_pp_it_1 ) : ( gb_pp_it_1 ) ;
assign n238 =  ( n27 ) ? ( gb_pp_it_1 ) : ( n237 ) ;
assign n239 =  ( n22 ) ? ( gb_pp_it_1 ) : ( n238 ) ;
assign n240 =  ( n13 ) ? ( 1'd1 ) : ( n239 ) ;
assign n241 =  ( n4 ) ? ( gb_pp_it_1 ) : ( n240 ) ;
assign n242 =  ( n38 ) ? ( gb_pp_it_2 ) : ( gb_pp_it_2 ) ;
assign n243 =  ( n27 ) ? ( gb_pp_it_2 ) : ( n242 ) ;
assign n244 =  ( n22 ) ? ( gb_pp_it_2 ) : ( n243 ) ;
assign n245 =  ( n13 ) ? ( gb_pp_it_1 ) : ( n244 ) ;
assign n246 =  ( n4 ) ? ( gb_pp_it_2 ) : ( n245 ) ;
assign n247 =  ( n38 ) ? ( gb_pp_it_3 ) : ( gb_pp_it_3 ) ;
assign n248 =  ( n27 ) ? ( gb_pp_it_3 ) : ( n247 ) ;
assign n249 =  ( n22 ) ? ( gb_pp_it_3 ) : ( n248 ) ;
assign n250 =  ( n13 ) ? ( gb_pp_it_2 ) : ( n249 ) ;
assign n251 =  ( n4 ) ? ( gb_pp_it_3 ) : ( n250 ) ;
assign n252 =  ( n38 ) ? ( gb_pp_it_4 ) : ( gb_pp_it_4 ) ;
assign n253 =  ( n27 ) ? ( gb_pp_it_4 ) : ( n252 ) ;
assign n254 =  ( n22 ) ? ( gb_pp_it_4 ) : ( n253 ) ;
assign n255 =  ( n13 ) ? ( gb_pp_it_3 ) : ( n254 ) ;
assign n256 =  ( n4 ) ? ( gb_pp_it_4 ) : ( n255 ) ;
assign n257 =  ( n38 ) ? ( gb_pp_it_5 ) : ( gb_pp_it_5 ) ;
assign n258 =  ( n27 ) ? ( gb_pp_it_5 ) : ( n257 ) ;
assign n259 =  ( n22 ) ? ( gb_pp_it_5 ) : ( n258 ) ;
assign n260 =  ( n13 ) ? ( gb_pp_it_4 ) : ( n259 ) ;
assign n261 =  ( n4 ) ? ( gb_pp_it_5 ) : ( n260 ) ;
assign n262 =  ( n38 ) ? ( gb_pp_it_6 ) : ( gb_pp_it_6 ) ;
assign n263 =  ( n27 ) ? ( gb_pp_it_6 ) : ( n262 ) ;
assign n264 =  ( n22 ) ? ( gb_pp_it_6 ) : ( n263 ) ;
assign n265 =  ( n13 ) ? ( gb_pp_it_5 ) : ( n264 ) ;
assign n266 =  ( n4 ) ? ( gb_pp_it_6 ) : ( n265 ) ;
assign n267 =  ( n38 ) ? ( gb_pp_it_7 ) : ( gb_pp_it_7 ) ;
assign n268 =  ( n27 ) ? ( gb_pp_it_7 ) : ( n267 ) ;
assign n269 =  ( n22 ) ? ( gb_pp_it_7 ) : ( n268 ) ;
assign n270 =  ( n13 ) ? ( gb_pp_it_6 ) : ( n269 ) ;
assign n271 =  ( n4 ) ? ( gb_pp_it_7 ) : ( n270 ) ;
assign n272 =  ( n38 ) ? ( gb_pp_it_8 ) : ( gb_pp_it_8 ) ;
assign n273 =  ( n27 ) ? ( gb_pp_it_8 ) : ( n272 ) ;
assign n274 =  ( n22 ) ? ( gb_pp_it_8 ) : ( n273 ) ;
assign n275 =  ( n13 ) ? ( gb_pp_it_7 ) : ( n274 ) ;
assign n276 =  ( n4 ) ? ( gb_pp_it_8 ) : ( n275 ) ;
assign n277 =  ( n38 ) ? ( gb_pp_it_9 ) : ( gb_pp_it_9 ) ;
assign n278 =  ( n27 ) ? ( gb_pp_it_9 ) : ( n277 ) ;
assign n279 =  ( n22 ) ? ( gb_pp_it_9 ) : ( n278 ) ;
assign n280 =  ( n13 ) ? ( gb_pp_it_8 ) : ( n279 ) ;
assign n281 =  ( n4 ) ? ( gb_pp_it_9 ) : ( n280 ) ;
assign n282 =  ( n38 ) ? ( LB1D_uIn ) : ( in_stream_buff_0 ) ;
assign n283 =  ( n33 ) ? ( LB1D_uIn ) : ( n282 ) ;
assign n284 =  ( n27 ) ? ( in_stream_buff_0 ) : ( n283 ) ;
assign n285 =  ( n22 ) ? ( in_stream_buff_0 ) : ( n284 ) ;
assign n286 =  ( n13 ) ? ( in_stream_buff_0 ) : ( n285 ) ;
assign n287 =  ( n4 ) ? ( in_stream_buff_0 ) : ( n286 ) ;
assign n288 =  ( n38 ) ? ( in_stream_buff_0 ) : ( in_stream_buff_1 ) ;
assign n289 =  ( n33 ) ? ( in_stream_buff_0 ) : ( n288 ) ;
assign n290 =  ( n27 ) ? ( in_stream_buff_1 ) : ( n289 ) ;
assign n291 =  ( n22 ) ? ( in_stream_buff_1 ) : ( n290 ) ;
assign n292 =  ( n13 ) ? ( in_stream_buff_1 ) : ( n291 ) ;
assign n293 =  ( n4 ) ? ( in_stream_buff_1 ) : ( n292 ) ;
assign n294 =  ( in_stream_full ) == ( 1'd1 )  ;
assign n295 =  ( n294 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n296 =  ( n38 ) ? ( 1'd0 ) : ( in_stream_empty ) ;
assign n297 =  ( n33 ) ? ( 1'd0 ) : ( n296 ) ;
assign n298 =  ( n27 ) ? ( n295 ) : ( n297 ) ;
assign n299 =  ( n22 ) ? ( in_stream_empty ) : ( n298 ) ;
assign n300 =  ( n13 ) ? ( in_stream_empty ) : ( n299 ) ;
assign n301 =  ( n4 ) ? ( in_stream_empty ) : ( n300 ) ;
assign n302 =  ( in_stream_empty ) == ( 1'd1 )  ;
assign n303 =  ( n302 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n304 =  ( n38 ) ? ( n303 ) : ( in_stream_full ) ;
assign n305 =  ( n33 ) ? ( n303 ) : ( n304 ) ;
assign n306 =  ( n27 ) ? ( 1'd0 ) : ( n305 ) ;
assign n307 =  ( n22 ) ? ( in_stream_full ) : ( n306 ) ;
assign n308 =  ( n13 ) ? ( in_stream_full ) : ( n307 ) ;
assign n309 =  ( n4 ) ? ( in_stream_full ) : ( n308 ) ;
assign n310 =  ( n294 ) ? ( in_stream_buff_1 ) : ( in_stream_buff_0 ) ;
assign n311 =  ( LB2D_proc_w ) == ( 64'd0 )  ;
assign n312 =  ( LB2D_proc_x ) - ( 9'd1 )  ;
assign n313 =  (  LB2D_proc_7 [ n312 ] )  ;
assign n314 =  ( LB2D_proc_w ) == ( 64'd1 )  ;
assign n315 =  (  LB2D_proc_0 [ n312 ] )  ;
assign n316 =  ( LB2D_proc_w ) == ( 64'd2 )  ;
assign n317 =  (  LB2D_proc_1 [ n312 ] )  ;
assign n318 =  ( LB2D_proc_w ) == ( 64'd3 )  ;
assign n319 =  (  LB2D_proc_2 [ n312 ] )  ;
assign n320 =  ( LB2D_proc_w ) == ( 64'd4 )  ;
assign n321 =  (  LB2D_proc_3 [ n312 ] )  ;
assign n322 =  ( LB2D_proc_w ) == ( 64'd5 )  ;
assign n323 =  (  LB2D_proc_4 [ n312 ] )  ;
assign n324 =  ( LB2D_proc_w ) == ( 64'd6 )  ;
assign n325 =  (  LB2D_proc_5 [ n312 ] )  ;
assign n326 =  (  LB2D_proc_6 [ n312 ] )  ;
assign n327 =  ( n324 ) ? ( n325 ) : ( n326 ) ;
assign n328 =  ( n322 ) ? ( n323 ) : ( n327 ) ;
assign n329 =  ( n320 ) ? ( n321 ) : ( n328 ) ;
assign n330 =  ( n318 ) ? ( n319 ) : ( n329 ) ;
assign n331 =  ( n316 ) ? ( n317 ) : ( n330 ) ;
assign n332 =  ( n314 ) ? ( n315 ) : ( n331 ) ;
assign n333 =  ( n311 ) ? ( n313 ) : ( n332 ) ;
assign n334 =  ( n324 ) ? ( n323 ) : ( n325 ) ;
assign n335 =  ( n322 ) ? ( n321 ) : ( n334 ) ;
assign n336 =  ( n320 ) ? ( n319 ) : ( n335 ) ;
assign n337 =  ( n318 ) ? ( n317 ) : ( n336 ) ;
assign n338 =  ( n316 ) ? ( n315 ) : ( n337 ) ;
assign n339 =  ( n314 ) ? ( n313 ) : ( n338 ) ;
assign n340 =  ( n311 ) ? ( n326 ) : ( n339 ) ;
assign n341 =  ( n324 ) ? ( n321 ) : ( n323 ) ;
assign n342 =  ( n322 ) ? ( n319 ) : ( n341 ) ;
assign n343 =  ( n320 ) ? ( n317 ) : ( n342 ) ;
assign n344 =  ( n318 ) ? ( n315 ) : ( n343 ) ;
assign n345 =  ( n316 ) ? ( n313 ) : ( n344 ) ;
assign n346 =  ( n314 ) ? ( n326 ) : ( n345 ) ;
assign n347 =  ( n311 ) ? ( n325 ) : ( n346 ) ;
assign n348 =  ( n324 ) ? ( n319 ) : ( n321 ) ;
assign n349 =  ( n322 ) ? ( n317 ) : ( n348 ) ;
assign n350 =  ( n320 ) ? ( n315 ) : ( n349 ) ;
assign n351 =  ( n318 ) ? ( n313 ) : ( n350 ) ;
assign n352 =  ( n316 ) ? ( n326 ) : ( n351 ) ;
assign n353 =  ( n314 ) ? ( n325 ) : ( n352 ) ;
assign n354 =  ( n311 ) ? ( n323 ) : ( n353 ) ;
assign n355 =  ( n324 ) ? ( n317 ) : ( n319 ) ;
assign n356 =  ( n322 ) ? ( n315 ) : ( n355 ) ;
assign n357 =  ( n320 ) ? ( n313 ) : ( n356 ) ;
assign n358 =  ( n318 ) ? ( n326 ) : ( n357 ) ;
assign n359 =  ( n316 ) ? ( n325 ) : ( n358 ) ;
assign n360 =  ( n314 ) ? ( n323 ) : ( n359 ) ;
assign n361 =  ( n311 ) ? ( n321 ) : ( n360 ) ;
assign n362 =  ( n324 ) ? ( n315 ) : ( n317 ) ;
assign n363 =  ( n322 ) ? ( n313 ) : ( n362 ) ;
assign n364 =  ( n320 ) ? ( n326 ) : ( n363 ) ;
assign n365 =  ( n318 ) ? ( n325 ) : ( n364 ) ;
assign n366 =  ( n316 ) ? ( n323 ) : ( n365 ) ;
assign n367 =  ( n314 ) ? ( n321 ) : ( n366 ) ;
assign n368 =  ( n311 ) ? ( n319 ) : ( n367 ) ;
assign n369 =  ( n324 ) ? ( n313 ) : ( n315 ) ;
assign n370 =  ( n322 ) ? ( n326 ) : ( n369 ) ;
assign n371 =  ( n320 ) ? ( n325 ) : ( n370 ) ;
assign n372 =  ( n318 ) ? ( n323 ) : ( n371 ) ;
assign n373 =  ( n316 ) ? ( n321 ) : ( n372 ) ;
assign n374 =  ( n314 ) ? ( n319 ) : ( n373 ) ;
assign n375 =  ( n311 ) ? ( n317 ) : ( n374 ) ;
assign n376 =  ( n324 ) ? ( n326 ) : ( n313 ) ;
assign n377 =  ( n322 ) ? ( n325 ) : ( n376 ) ;
assign n378 =  ( n320 ) ? ( n323 ) : ( n377 ) ;
assign n379 =  ( n318 ) ? ( n321 ) : ( n378 ) ;
assign n380 =  ( n316 ) ? ( n319 ) : ( n379 ) ;
assign n381 =  ( n314 ) ? ( n317 ) : ( n380 ) ;
assign n382 =  ( n311 ) ? ( n315 ) : ( n381 ) ;
assign n383 =  { ( n375 ) , ( n382 ) }  ;
assign n384 =  { ( n368 ) , ( n383 ) }  ;
assign n385 =  { ( n361 ) , ( n384 ) }  ;
assign n386 =  { ( n354 ) , ( n385 ) }  ;
assign n387 =  { ( n347 ) , ( n386 ) }  ;
assign n388 =  { ( n340 ) , ( n387 ) }  ;
assign n389 =  { ( n333 ) , ( n388 ) }  ;
assign n390 =  { ( n310 ) , ( n389 ) }  ;
assign n391 =  ( n25 ) ? ( slice_stream_buff_0 ) : ( n390 ) ;
assign n392 =  ( n38 ) ? ( slice_stream_buff_0 ) : ( slice_stream_buff_0 ) ;
assign n393 =  ( n27 ) ? ( n391 ) : ( n392 ) ;
assign n394 =  ( n22 ) ? ( slice_stream_buff_0 ) : ( n393 ) ;
assign n395 =  ( n13 ) ? ( slice_stream_buff_0 ) : ( n394 ) ;
assign n396 =  ( n4 ) ? ( slice_stream_buff_0 ) : ( n395 ) ;
assign n397 =  ( n25 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n398 =  ( n38 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_1 ) ;
assign n399 =  ( n27 ) ? ( n397 ) : ( n398 ) ;
assign n400 =  ( n22 ) ? ( slice_stream_buff_1 ) : ( n399 ) ;
assign n401 =  ( n13 ) ? ( slice_stream_buff_1 ) : ( n400 ) ;
assign n402 =  ( n4 ) ? ( slice_stream_buff_1 ) : ( n401 ) ;
assign n403 =  ( n135 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n404 =  ( n25 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n405 =  ( n38 ) ? ( slice_stream_empty ) : ( slice_stream_empty ) ;
assign n406 =  ( n27 ) ? ( n404 ) : ( n405 ) ;
assign n407 =  ( n22 ) ? ( n403 ) : ( n406 ) ;
assign n408 =  ( n13 ) ? ( slice_stream_empty ) : ( n407 ) ;
assign n409 =  ( n4 ) ? ( slice_stream_empty ) : ( n408 ) ;
assign n410 =  ( slice_stream_empty ) == ( 1'd1 )  ;
assign n411 =  ( n410 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n412 =  ( n25 ) ? ( 1'd0 ) : ( n411 ) ;
assign n413 =  ( n38 ) ? ( slice_stream_full ) : ( slice_stream_full ) ;
assign n414 =  ( n27 ) ? ( n412 ) : ( n413 ) ;
assign n415 =  ( n22 ) ? ( 1'd0 ) : ( n414 ) ;
assign n416 =  ( n13 ) ? ( slice_stream_full ) : ( n415 ) ;
assign n417 =  ( n4 ) ? ( slice_stream_full ) : ( n416 ) ;
assign n418 =  ( LB2D_shift_x ) >= ( 9'd8 )  ;
assign n419 =  ( LB2D_shift_x ) == ( 9'd0 )  ;
assign n420 =  ( n418 ) | ( n419 )  ;
assign n421 = n136[71:64] ;
assign n422 = LB2D_shift_7[71:64] ;
assign n423 = LB2D_shift_6[71:64] ;
assign n424 = LB2D_shift_5[71:64] ;
assign n425 = LB2D_shift_4[71:64] ;
assign n426 = LB2D_shift_3[71:64] ;
assign n427 = LB2D_shift_2[71:64] ;
assign n428 = LB2D_shift_1[71:64] ;
assign n429 = LB2D_shift_0[71:64] ;
assign n430 =  { ( n428 ) , ( n429 ) }  ;
assign n431 =  { ( n427 ) , ( n430 ) }  ;
assign n432 =  { ( n426 ) , ( n431 ) }  ;
assign n433 =  { ( n425 ) , ( n432 ) }  ;
assign n434 =  { ( n424 ) , ( n433 ) }  ;
assign n435 =  { ( n423 ) , ( n434 ) }  ;
assign n436 =  { ( n422 ) , ( n435 ) }  ;
assign n437 =  { ( n421 ) , ( n436 ) }  ;
assign n438 = n136[63:56] ;
assign n439 = LB2D_shift_7[63:56] ;
assign n440 = LB2D_shift_6[63:56] ;
assign n441 = LB2D_shift_5[63:56] ;
assign n442 = LB2D_shift_4[63:56] ;
assign n443 = LB2D_shift_3[63:56] ;
assign n444 = LB2D_shift_2[63:56] ;
assign n445 = LB2D_shift_1[63:56] ;
assign n446 = LB2D_shift_0[63:56] ;
assign n447 =  { ( n445 ) , ( n446 ) }  ;
assign n448 =  { ( n444 ) , ( n447 ) }  ;
assign n449 =  { ( n443 ) , ( n448 ) }  ;
assign n450 =  { ( n442 ) , ( n449 ) }  ;
assign n451 =  { ( n441 ) , ( n450 ) }  ;
assign n452 =  { ( n440 ) , ( n451 ) }  ;
assign n453 =  { ( n439 ) , ( n452 ) }  ;
assign n454 =  { ( n438 ) , ( n453 ) }  ;
assign n455 = n136[55:48] ;
assign n456 = LB2D_shift_7[55:48] ;
assign n457 = LB2D_shift_6[55:48] ;
assign n458 = LB2D_shift_5[55:48] ;
assign n459 = LB2D_shift_4[55:48] ;
assign n460 = LB2D_shift_3[55:48] ;
assign n461 = LB2D_shift_2[55:48] ;
assign n462 = LB2D_shift_1[55:48] ;
assign n463 = LB2D_shift_0[55:48] ;
assign n464 =  { ( n462 ) , ( n463 ) }  ;
assign n465 =  { ( n461 ) , ( n464 ) }  ;
assign n466 =  { ( n460 ) , ( n465 ) }  ;
assign n467 =  { ( n459 ) , ( n466 ) }  ;
assign n468 =  { ( n458 ) , ( n467 ) }  ;
assign n469 =  { ( n457 ) , ( n468 ) }  ;
assign n470 =  { ( n456 ) , ( n469 ) }  ;
assign n471 =  { ( n455 ) , ( n470 ) }  ;
assign n472 = n136[47:40] ;
assign n473 = LB2D_shift_7[47:40] ;
assign n474 = LB2D_shift_6[47:40] ;
assign n475 = LB2D_shift_5[47:40] ;
assign n476 = LB2D_shift_4[47:40] ;
assign n477 = LB2D_shift_3[47:40] ;
assign n478 = LB2D_shift_2[47:40] ;
assign n479 = LB2D_shift_1[47:40] ;
assign n480 = LB2D_shift_0[47:40] ;
assign n481 =  { ( n479 ) , ( n480 ) }  ;
assign n482 =  { ( n478 ) , ( n481 ) }  ;
assign n483 =  { ( n477 ) , ( n482 ) }  ;
assign n484 =  { ( n476 ) , ( n483 ) }  ;
assign n485 =  { ( n475 ) , ( n484 ) }  ;
assign n486 =  { ( n474 ) , ( n485 ) }  ;
assign n487 =  { ( n473 ) , ( n486 ) }  ;
assign n488 =  { ( n472 ) , ( n487 ) }  ;
assign n489 = n136[39:32] ;
assign n490 = LB2D_shift_7[39:32] ;
assign n491 = LB2D_shift_6[39:32] ;
assign n492 = LB2D_shift_5[39:32] ;
assign n493 = LB2D_shift_4[39:32] ;
assign n494 = LB2D_shift_3[39:32] ;
assign n495 = LB2D_shift_2[39:32] ;
assign n496 = LB2D_shift_1[39:32] ;
assign n497 = LB2D_shift_0[39:32] ;
assign n498 =  { ( n496 ) , ( n497 ) }  ;
assign n499 =  { ( n495 ) , ( n498 ) }  ;
assign n500 =  { ( n494 ) , ( n499 ) }  ;
assign n501 =  { ( n493 ) , ( n500 ) }  ;
assign n502 =  { ( n492 ) , ( n501 ) }  ;
assign n503 =  { ( n491 ) , ( n502 ) }  ;
assign n504 =  { ( n490 ) , ( n503 ) }  ;
assign n505 =  { ( n489 ) , ( n504 ) }  ;
assign n506 = n136[31:24] ;
assign n507 = LB2D_shift_7[31:24] ;
assign n508 = LB2D_shift_6[31:24] ;
assign n509 = LB2D_shift_5[31:24] ;
assign n510 = LB2D_shift_4[31:24] ;
assign n511 = LB2D_shift_3[31:24] ;
assign n512 = LB2D_shift_2[31:24] ;
assign n513 = LB2D_shift_1[31:24] ;
assign n514 = LB2D_shift_0[31:24] ;
assign n515 =  { ( n513 ) , ( n514 ) }  ;
assign n516 =  { ( n512 ) , ( n515 ) }  ;
assign n517 =  { ( n511 ) , ( n516 ) }  ;
assign n518 =  { ( n510 ) , ( n517 ) }  ;
assign n519 =  { ( n509 ) , ( n518 ) }  ;
assign n520 =  { ( n508 ) , ( n519 ) }  ;
assign n521 =  { ( n507 ) , ( n520 ) }  ;
assign n522 =  { ( n506 ) , ( n521 ) }  ;
assign n523 = n136[23:16] ;
assign n524 = LB2D_shift_7[23:16] ;
assign n525 = LB2D_shift_6[23:16] ;
assign n526 = LB2D_shift_5[23:16] ;
assign n527 = LB2D_shift_4[23:16] ;
assign n528 = LB2D_shift_3[23:16] ;
assign n529 = LB2D_shift_2[23:16] ;
assign n530 = LB2D_shift_1[23:16] ;
assign n531 = LB2D_shift_0[23:16] ;
assign n532 =  { ( n530 ) , ( n531 ) }  ;
assign n533 =  { ( n529 ) , ( n532 ) }  ;
assign n534 =  { ( n528 ) , ( n533 ) }  ;
assign n535 =  { ( n527 ) , ( n534 ) }  ;
assign n536 =  { ( n526 ) , ( n535 ) }  ;
assign n537 =  { ( n525 ) , ( n536 ) }  ;
assign n538 =  { ( n524 ) , ( n537 ) }  ;
assign n539 =  { ( n523 ) , ( n538 ) }  ;
assign n540 = n136[15:8] ;
assign n541 = LB2D_shift_7[15:8] ;
assign n542 = LB2D_shift_6[15:8] ;
assign n543 = LB2D_shift_5[15:8] ;
assign n544 = LB2D_shift_4[15:8] ;
assign n545 = LB2D_shift_3[15:8] ;
assign n546 = LB2D_shift_2[15:8] ;
assign n547 = LB2D_shift_1[15:8] ;
assign n548 = LB2D_shift_0[15:8] ;
assign n549 =  { ( n547 ) , ( n548 ) }  ;
assign n550 =  { ( n546 ) , ( n549 ) }  ;
assign n551 =  { ( n545 ) , ( n550 ) }  ;
assign n552 =  { ( n544 ) , ( n551 ) }  ;
assign n553 =  { ( n543 ) , ( n552 ) }  ;
assign n554 =  { ( n542 ) , ( n553 ) }  ;
assign n555 =  { ( n541 ) , ( n554 ) }  ;
assign n556 =  { ( n540 ) , ( n555 ) }  ;
assign n557 = n136[7:0] ;
assign n558 = LB2D_shift_7[7:0] ;
assign n559 = LB2D_shift_6[7:0] ;
assign n560 = LB2D_shift_5[7:0] ;
assign n561 = LB2D_shift_4[7:0] ;
assign n562 = LB2D_shift_3[7:0] ;
assign n563 = LB2D_shift_2[7:0] ;
assign n564 = LB2D_shift_1[7:0] ;
assign n565 = LB2D_shift_0[7:0] ;
assign n566 =  { ( n564 ) , ( n565 ) }  ;
assign n567 =  { ( n563 ) , ( n566 ) }  ;
assign n568 =  { ( n562 ) , ( n567 ) }  ;
assign n569 =  { ( n561 ) , ( n568 ) }  ;
assign n570 =  { ( n560 ) , ( n569 ) }  ;
assign n571 =  { ( n559 ) , ( n570 ) }  ;
assign n572 =  { ( n558 ) , ( n571 ) }  ;
assign n573 =  { ( n557 ) , ( n572 ) }  ;
assign n574 =  { ( n556 ) , ( n573 ) }  ;
assign n575 =  { ( n539 ) , ( n574 ) }  ;
assign n576 =  { ( n522 ) , ( n575 ) }  ;
assign n577 =  { ( n505 ) , ( n576 ) }  ;
assign n578 =  { ( n488 ) , ( n577 ) }  ;
assign n579 =  { ( n471 ) , ( n578 ) }  ;
assign n580 =  { ( n454 ) , ( n579 ) }  ;
assign n581 =  { ( n437 ) , ( n580 ) }  ;
assign n582 =  ( n420 ) ? ( n581 ) : ( stencil_stream_buff_0 ) ;
assign n583 =  ( n38 ) ? ( stencil_stream_buff_0 ) : ( stencil_stream_buff_0 ) ;
assign n584 =  ( n27 ) ? ( stencil_stream_buff_0 ) : ( n583 ) ;
assign n585 =  ( n22 ) ? ( n582 ) : ( n584 ) ;
assign n586 =  ( n13 ) ? ( stencil_stream_buff_0 ) : ( n585 ) ;
assign n587 =  ( n4 ) ? ( stencil_stream_buff_0 ) : ( n586 ) ;
assign n588 =  ( n38 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_1 ) ;
assign n589 =  ( n27 ) ? ( stencil_stream_buff_1 ) : ( n588 ) ;
assign n590 =  ( n22 ) ? ( stencil_stream_buff_0 ) : ( n589 ) ;
assign n591 =  ( n13 ) ? ( stencil_stream_buff_1 ) : ( n590 ) ;
assign n592 =  ( n4 ) ? ( stencil_stream_buff_1 ) : ( n591 ) ;
assign n593 =  ( n163 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n594 = ~ ( n420 ) ;
assign n595 =  ( n594 ) ? ( stencil_stream_empty ) : ( 1'd0 ) ;
assign n596 =  ( n38 ) ? ( stencil_stream_empty ) : ( stencil_stream_empty ) ;
assign n597 =  ( n27 ) ? ( stencil_stream_empty ) : ( n596 ) ;
assign n598 =  ( n22 ) ? ( n595 ) : ( n597 ) ;
assign n599 =  ( n13 ) ? ( n593 ) : ( n598 ) ;
assign n600 =  ( n4 ) ? ( stencil_stream_empty ) : ( n599 ) ;
assign n601 =  ( n9 ) ? ( 1'd0 ) : ( 1'd0 ) ;
assign n602 =  ( stencil_stream_empty ) == ( 1'd1 )  ;
assign n603 =  ( n602 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n604 =  ( n594 ) ? ( stencil_stream_full ) : ( n603 ) ;
assign n605 =  ( n38 ) ? ( stencil_stream_full ) : ( stencil_stream_full ) ;
assign n606 =  ( n27 ) ? ( stencil_stream_full ) : ( n605 ) ;
assign n607 =  ( n22 ) ? ( n604 ) : ( n606 ) ;
assign n608 =  ( n13 ) ? ( n601 ) : ( n607 ) ;
assign n609 =  ( n4 ) ? ( stencil_stream_full ) : ( n608 ) ;
assign n610 = ~ ( n4 ) ;
assign n611 = ~ ( n13 ) ;
assign n612 =  ( n610 ) & ( n611 )  ;
assign n613 = ~ ( n22 ) ;
assign n614 =  ( n612 ) & ( n613 )  ;
assign n615 = ~ ( n27 ) ;
assign n616 =  ( n614 ) & ( n615 )  ;
assign n617 = ~ ( n38 ) ;
assign n618 =  ( n616 ) & ( n617 )  ;
assign n619 =  ( n616 ) & ( n38 )  ;
assign n620 =  ( n614 ) & ( n27 )  ;
assign n621 = ~ ( n311 ) ;
assign n622 =  ( n620 ) & ( n621 )  ;
assign n623 =  ( n620 ) & ( n311 )  ;
assign n624 =  ( n612 ) & ( n22 )  ;
assign n625 =  ( n610 ) & ( n13 )  ;
assign LB2D_proc_0_addr0 = n623 ? (n312) : (0);
assign LB2D_proc_0_data0 = n623 ? (n310) : (LB2D_proc_0[0]);
assign n626 = ~ ( n314 ) ;
assign n627 =  ( n620 ) & ( n626 )  ;
assign n628 =  ( n620 ) & ( n314 )  ;
assign LB2D_proc_1_addr0 = n628 ? (n312) : (0);
assign LB2D_proc_1_data0 = n628 ? (n310) : (LB2D_proc_1[0]);
assign n629 = ~ ( n316 ) ;
assign n630 =  ( n620 ) & ( n629 )  ;
assign n631 =  ( n620 ) & ( n316 )  ;
assign LB2D_proc_2_addr0 = n631 ? (n312) : (0);
assign LB2D_proc_2_data0 = n631 ? (n310) : (LB2D_proc_2[0]);
assign n632 = ~ ( n318 ) ;
assign n633 =  ( n620 ) & ( n632 )  ;
assign n634 =  ( n620 ) & ( n318 )  ;
assign LB2D_proc_3_addr0 = n634 ? (n312) : (0);
assign LB2D_proc_3_data0 = n634 ? (n310) : (LB2D_proc_3[0]);
assign n635 = ~ ( n320 ) ;
assign n636 =  ( n620 ) & ( n635 )  ;
assign n637 =  ( n620 ) & ( n320 )  ;
assign LB2D_proc_4_addr0 = n637 ? (n312) : (0);
assign LB2D_proc_4_data0 = n637 ? (n310) : (LB2D_proc_4[0]);
assign n638 = ~ ( n322 ) ;
assign n639 =  ( n620 ) & ( n638 )  ;
assign n640 =  ( n620 ) & ( n322 )  ;
assign LB2D_proc_5_addr0 = n640 ? (n312) : (0);
assign LB2D_proc_5_data0 = n640 ? (n310) : (LB2D_proc_5[0]);
assign n641 = ~ ( n324 ) ;
assign n642 =  ( n620 ) & ( n641 )  ;
assign n643 =  ( n620 ) & ( n324 )  ;
assign LB2D_proc_6_addr0 = n643 ? (n312) : (0);
assign LB2D_proc_6_data0 = n643 ? (n310) : (LB2D_proc_6[0]);
assign n644 = ~ ( n75 ) ;
assign n645 =  ( n620 ) & ( n644 )  ;
assign n646 =  ( n620 ) & ( n75 )  ;
assign LB2D_proc_7_addr0 = n646 ? (n312) : (0);
assign LB2D_proc_7_data0 = n646 ? (n310) : (LB2D_proc_7[0]);
/*
function [7:0] gb_fun ;
input [647:0] arg0;
    begin
//TODO: Add the specific function HERE.    end
endfunction
*/

always @(posedge clk) begin
   if(rst) begin
       LB1D_buff <= LB1D_buff;
       LB1D_in <= LB1D_in;
       LB1D_it_1 <= LB1D_it_1;
       LB1D_p_cnt <= LB1D_p_cnt;
       LB1D_uIn <= LB1D_uIn;
       LB2D_proc_w <= LB2D_proc_w;
       LB2D_proc_x <= LB2D_proc_x;
       LB2D_proc_y <= LB2D_proc_y;
       LB2D_shift_0 <= LB2D_shift_0;
       LB2D_shift_1 <= LB2D_shift_1;
       LB2D_shift_2 <= LB2D_shift_2;
       LB2D_shift_3 <= LB2D_shift_3;
       LB2D_shift_4 <= LB2D_shift_4;
       LB2D_shift_5 <= LB2D_shift_5;
       LB2D_shift_6 <= LB2D_shift_6;
       LB2D_shift_7 <= LB2D_shift_7;
       LB2D_shift_x <= LB2D_shift_x;
       LB2D_shift_y <= LB2D_shift_y;
       arg_0_TDATA <= arg_0_TDATA;
       arg_0_TVALID <= arg_0_TVALID;
       arg_1_TREADY <= arg_1_TREADY;
       gb_exit_it_1 <= gb_exit_it_1;
       gb_exit_it_2 <= gb_exit_it_2;
       gb_exit_it_3 <= gb_exit_it_3;
       gb_exit_it_4 <= gb_exit_it_4;
       gb_exit_it_5 <= gb_exit_it_5;
       gb_exit_it_6 <= gb_exit_it_6;
       gb_exit_it_7 <= gb_exit_it_7;
       gb_exit_it_8 <= gb_exit_it_8;
       gb_p_cnt <= gb_p_cnt;
       gb_pp_it_1 <= gb_pp_it_1;
       gb_pp_it_2 <= gb_pp_it_2;
       gb_pp_it_3 <= gb_pp_it_3;
       gb_pp_it_4 <= gb_pp_it_4;
       gb_pp_it_5 <= gb_pp_it_5;
       gb_pp_it_6 <= gb_pp_it_6;
       gb_pp_it_7 <= gb_pp_it_7;
       gb_pp_it_8 <= gb_pp_it_8;
       gb_pp_it_9 <= gb_pp_it_9;
       in_stream_buff_0 <= in_stream_buff_0;
       in_stream_buff_1 <= in_stream_buff_1;
       in_stream_empty <= in_stream_empty;
       in_stream_full <= in_stream_full;
       slice_stream_buff_0 <= slice_stream_buff_0;
       slice_stream_buff_1 <= slice_stream_buff_1;
       slice_stream_empty <= slice_stream_empty;
       slice_stream_full <= slice_stream_full;
       stencil_stream_buff_0 <= stencil_stream_buff_0;
       stencil_stream_buff_1 <= stencil_stream_buff_1;
       stencil_stream_empty <= stencil_stream_empty;
       stencil_stream_full <= stencil_stream_full;
   end
   else if(step) begin
       LB1D_buff <= n45;
       LB1D_in <= n52;
       LB1D_it_1 <= n58;
       LB1D_p_cnt <= n66;
       LB1D_uIn <= n73;
       LB2D_proc_w <= n83;
       LB2D_proc_x <= n90;
       LB2D_proc_y <= n99;
       LB2D_shift_0 <= n104;
       LB2D_shift_1 <= n109;
       LB2D_shift_2 <= n114;
       LB2D_shift_3 <= n119;
       LB2D_shift_4 <= n124;
       LB2D_shift_5 <= n129;
       LB2D_shift_6 <= n134;
       LB2D_shift_7 <= n141;
       LB2D_shift_x <= n152;
       LB2D_shift_y <= n162;
       arg_0_TDATA <= n171;
       arg_0_TVALID <= n179;
       arg_1_TREADY <= n186;
       gb_exit_it_1 <= n194;
       gb_exit_it_2 <= n199;
       gb_exit_it_3 <= n204;
       gb_exit_it_4 <= n209;
       gb_exit_it_5 <= n214;
       gb_exit_it_6 <= n219;
       gb_exit_it_7 <= n224;
       gb_exit_it_8 <= n229;
       gb_p_cnt <= n236;
       gb_pp_it_1 <= n241;
       gb_pp_it_2 <= n246;
       gb_pp_it_3 <= n251;
       gb_pp_it_4 <= n256;
       gb_pp_it_5 <= n261;
       gb_pp_it_6 <= n266;
       gb_pp_it_7 <= n271;
       gb_pp_it_8 <= n276;
       gb_pp_it_9 <= n281;
       in_stream_buff_0 <= n287;
       in_stream_buff_1 <= n293;
       in_stream_empty <= n301;
       in_stream_full <= n309;
       slice_stream_buff_0 <= n396;
       slice_stream_buff_1 <= n402;
       slice_stream_empty <= n409;
       slice_stream_full <= n417;
       stencil_stream_buff_0 <= n587;
       stencil_stream_buff_1 <= n592;
       stencil_stream_empty <= n600;
       stencil_stream_full <= n609;
       LB2D_proc_0 [ LB2D_proc_0_addr0 ] <= LB2D_proc_0_data0;
       LB2D_proc_1 [ LB2D_proc_1_addr0 ] <= LB2D_proc_1_data0;
       LB2D_proc_2 [ LB2D_proc_2_addr0 ] <= LB2D_proc_2_data0;
       LB2D_proc_3 [ LB2D_proc_3_addr0 ] <= LB2D_proc_3_data0;
       LB2D_proc_4 [ LB2D_proc_4_addr0 ] <= LB2D_proc_4_data0;
       LB2D_proc_5 [ LB2D_proc_5_addr0 ] <= LB2D_proc_5_data0;
       LB2D_proc_6 [ LB2D_proc_6_addr0 ] <= LB2D_proc_6_data0;
       LB2D_proc_7 [ LB2D_proc_7_addr0 ] <= LB2D_proc_7_data0;
   end
end
endmodule
