module SPEC_B(
arg_0_TREADY,
arg_1_TDATA,
arg_1_TVALID,
LB1D_buff,
LB1D_in,
LB1D_it_1,
LB1D_p_cnt,
LB1D_uIn,
LB2D_proc_w,
LB2D_proc_x,
LB2D_proc_y,
LB2D_shift_0,
LB2D_shift_1,
LB2D_shift_2,
LB2D_shift_3,
LB2D_shift_4,
LB2D_shift_5,
LB2D_shift_6,
LB2D_shift_7,
LB2D_shift_x,
LB2D_shift_y,
arg_0_TDATA,
arg_0_TVALID,
arg_1_TREADY,
gb_exit_it_1,
gb_exit_it_2,
gb_exit_it_3,
gb_exit_it_4,
gb_exit_it_5,
gb_exit_it_6,
gb_exit_it_7,
gb_exit_it_8,
gb_p_cnt,
gb_pp_it_1,
gb_pp_it_2,
gb_pp_it_3,
gb_pp_it_4,
gb_pp_it_5,
gb_pp_it_6,
gb_pp_it_7,
gb_pp_it_8,
gb_pp_it_9,
in_stream_buff_0,
in_stream_buff_1,
in_stream_empty,
in_stream_full,
slice_stream_buff_0,
slice_stream_buff_1,
slice_stream_empty,
slice_stream_full,
stencil_stream_buff_0,
stencil_stream_buff_1,
stencil_stream_empty,
stencil_stream_full,
clk,rst,
step
);
input            arg_0_TREADY;
input      [7:0] arg_1_TDATA;
input            arg_1_TVALID;
input clk;
input rst;
input step;
output      [7:0] LB1D_buff;
output      [7:0] LB1D_in;
output            LB1D_it_1;
output     [18:0] LB1D_p_cnt;
output      [7:0] LB1D_uIn;
output     [63:0] LB2D_proc_w;
output      [8:0] LB2D_proc_x;
output      [9:0] LB2D_proc_y;
output     [71:0] LB2D_shift_0;
output     [71:0] LB2D_shift_1;
output     [71:0] LB2D_shift_2;
output     [71:0] LB2D_shift_3;
output     [71:0] LB2D_shift_4;
output     [71:0] LB2D_shift_5;
output     [71:0] LB2D_shift_6;
output     [71:0] LB2D_shift_7;
output      [8:0] LB2D_shift_x;
output      [9:0] LB2D_shift_y;
output      [7:0] arg_0_TDATA;
output            arg_0_TVALID;
output            arg_1_TREADY;
output            gb_exit_it_1;
output            gb_exit_it_2;
output            gb_exit_it_3;
output            gb_exit_it_4;
output            gb_exit_it_5;
output            gb_exit_it_6;
output            gb_exit_it_7;
output            gb_exit_it_8;
output     [18:0] gb_p_cnt;
output            gb_pp_it_1;
output            gb_pp_it_2;
output            gb_pp_it_3;
output            gb_pp_it_4;
output            gb_pp_it_5;
output            gb_pp_it_6;
output            gb_pp_it_7;
output            gb_pp_it_8;
output            gb_pp_it_9;
output      [7:0] in_stream_buff_0;
output      [7:0] in_stream_buff_1;
output            in_stream_empty;
output            in_stream_full;
output     [71:0] slice_stream_buff_0;
output     [71:0] slice_stream_buff_1;
output            slice_stream_empty;
output            slice_stream_full;
output    [647:0] stencil_stream_buff_0;
output    [647:0] stencil_stream_buff_1;
output            stencil_stream_empty;
output            stencil_stream_full;
reg      [7:0] LB1D_buff;
reg      [7:0] LB1D_in;
reg            LB1D_it_1;
reg     [18:0] LB1D_p_cnt;
reg      [7:0] LB1D_uIn;
reg     [63:0] LB2D_proc_w;
reg      [8:0] LB2D_proc_x;
reg      [9:0] LB2D_proc_y;
reg     [71:0] LB2D_shift_0;
reg     [71:0] LB2D_shift_1;
reg     [71:0] LB2D_shift_2;
reg     [71:0] LB2D_shift_3;
reg     [71:0] LB2D_shift_4;
reg     [71:0] LB2D_shift_5;
reg     [71:0] LB2D_shift_6;
reg     [71:0] LB2D_shift_7;
reg      [8:0] LB2D_shift_x;
reg      [9:0] LB2D_shift_y;
reg      [7:0] arg_0_TDATA;
reg            arg_0_TVALID;
reg            arg_1_TREADY;
reg            gb_exit_it_1;
reg            gb_exit_it_2;
reg            gb_exit_it_3;
reg            gb_exit_it_4;
reg            gb_exit_it_5;
reg            gb_exit_it_6;
reg            gb_exit_it_7;
reg            gb_exit_it_8;
reg     [18:0] gb_p_cnt;
reg            gb_pp_it_1;
reg            gb_pp_it_2;
reg            gb_pp_it_3;
reg            gb_pp_it_4;
reg            gb_pp_it_5;
reg            gb_pp_it_6;
reg            gb_pp_it_7;
reg            gb_pp_it_8;
reg            gb_pp_it_9;
reg      [7:0] in_stream_buff_0;
reg      [7:0] in_stream_buff_1;
reg            in_stream_empty;
reg            in_stream_full;
reg     [71:0] slice_stream_buff_0;
reg     [71:0] slice_stream_buff_1;
reg            slice_stream_empty;
reg            slice_stream_full;
reg    [647:0] stencil_stream_buff_0;
reg    [647:0] stencil_stream_buff_1;
reg            stencil_stream_empty;
reg            stencil_stream_full;
wire            arg_0_TREADY;
wire      [7:0] arg_1_TDATA;
wire            arg_1_TVALID;
wire            n0;
wire            n1;
wire            n2;
wire            n3;
wire            n4;
wire            n5;
wire            n6;
wire            n7;
wire            n8;
wire            n9;
wire            n10;
wire            n11;
wire            n12;
wire            n13;
wire            n14;
wire            n15;
wire            n16;
wire            n17;
wire            n18;
wire            n19;
wire            n20;
wire            n21;
wire            n22;
wire            n23;
wire            n24;
wire            n25;
wire            n26;
wire            n27;
wire            n28;
wire            n29;
wire            n30;
wire            n31;
wire            n32;
wire      [7:0] n33;
wire      [7:0] n34;
wire      [7:0] n35;
wire      [7:0] n36;
wire      [7:0] n37;
wire      [7:0] n38;
wire      [7:0] n39;
wire      [7:0] n40;
wire      [7:0] n41;
wire      [7:0] n42;
wire      [7:0] n43;
wire      [7:0] n44;
wire            n45;
wire     [18:0] n46;
wire     [18:0] n47;
wire            n48;
wire     [18:0] n49;
wire     [18:0] n50;
wire     [18:0] n51;
wire     [18:0] n52;
wire     [18:0] n53;
wire     [18:0] n54;
wire     [18:0] n55;
wire      [7:0] n56;
wire      [7:0] n57;
wire      [7:0] n58;
wire      [7:0] n59;
wire      [7:0] n60;
wire      [7:0] n61;
wire            n62;
wire            n63;
wire     [63:0] n64;
wire     [63:0] n65;
wire     [63:0] n66;
wire     [63:0] n67;
wire     [63:0] n68;
wire     [63:0] n69;
wire     [63:0] n70;
wire     [63:0] n71;
wire      [8:0] n72;
wire      [8:0] n73;
wire      [8:0] n74;
wire      [8:0] n75;
wire      [8:0] n76;
wire      [8:0] n77;
wire      [8:0] n78;
wire            n79;
wire      [9:0] n80;
wire      [9:0] n81;
wire      [9:0] n82;
wire      [9:0] n83;
wire      [9:0] n84;
wire      [9:0] n85;
wire      [9:0] n86;
wire      [9:0] n87;
wire     [71:0] n88;
wire     [71:0] n89;
wire     [71:0] n90;
wire     [71:0] n91;
wire     [71:0] n92;
wire     [71:0] n93;
wire     [71:0] n94;
wire     [71:0] n95;
wire     [71:0] n96;
wire     [71:0] n97;
wire     [71:0] n98;
wire     [71:0] n99;
wire     [71:0] n100;
wire     [71:0] n101;
wire     [71:0] n102;
wire     [71:0] n103;
wire     [71:0] n104;
wire     [71:0] n105;
wire     [71:0] n106;
wire     [71:0] n107;
wire     [71:0] n108;
wire     [71:0] n109;
wire     [71:0] n110;
wire     [71:0] n111;
wire     [71:0] n112;
wire     [71:0] n113;
wire     [71:0] n114;
wire     [71:0] n115;
wire     [71:0] n116;
wire     [71:0] n117;
wire     [71:0] n118;
wire     [71:0] n119;
wire     [71:0] n120;
wire     [71:0] n121;
wire     [71:0] n122;
wire            n123;
wire     [71:0] n124;
wire     [71:0] n125;
wire     [71:0] n126;
wire     [71:0] n127;
wire     [71:0] n128;
wire     [71:0] n129;
wire            n130;
wire            n131;
wire            n132;
wire      [8:0] n133;
wire      [8:0] n134;
wire      [8:0] n135;
wire      [8:0] n136;
wire      [8:0] n137;
wire      [8:0] n138;
wire      [8:0] n139;
wire            n140;
wire            n141;
wire      [9:0] n142;
wire      [9:0] n143;
wire      [9:0] n144;
wire      [9:0] n145;
wire      [9:0] n146;
wire      [9:0] n147;
wire      [9:0] n148;
wire      [9:0] n149;
wire            n150;
wire    [647:0] n151;
wire      [7:0] n152;
wire      [7:0] n153;
wire      [7:0] n154;
wire      [7:0] n155;
wire      [7:0] n156;
wire      [7:0] n157;
wire            n158;
wire            n159;
wire            n160;
wire            n161;
wire            n162;
wire            n163;
wire            n164;
wire            n165;
wire            n166;
wire            n167;
wire            n168;
wire            n169;
wire            n170;
wire     [18:0] n171;
wire            n172;
wire            n173;
wire            n174;
wire            n175;
wire            n176;
wire            n177;
wire            n178;
wire            n179;
wire            n180;
wire            n181;
wire            n182;
wire            n183;
wire            n184;
wire            n185;
wire            n186;
wire            n187;
wire            n188;
wire            n189;
wire            n190;
wire            n191;
wire            n192;
wire            n193;
wire            n194;
wire            n195;
wire            n196;
wire            n197;
wire            n198;
wire            n199;
wire            n200;
wire            n201;
wire            n202;
wire            n203;
wire            n204;
wire            n205;
wire            n206;
wire            n207;
wire            n208;
wire            n209;
wire            n210;
wire            n211;
wire            n212;
wire            n213;
wire            n214;
wire     [18:0] n215;
wire     [18:0] n216;
wire     [18:0] n217;
wire     [18:0] n218;
wire     [18:0] n219;
wire     [18:0] n220;
wire            n221;
wire            n222;
wire            n223;
wire            n224;
wire            n225;
wire            n226;
wire            n227;
wire            n228;
wire            n229;
wire            n230;
wire            n231;
wire            n232;
wire            n233;
wire            n234;
wire            n235;
wire            n236;
wire            n237;
wire            n238;
wire            n239;
wire            n240;
wire            n241;
wire            n242;
wire            n243;
wire            n244;
wire            n245;
wire            n246;
wire            n247;
wire            n248;
wire            n249;
wire            n250;
wire            n251;
wire            n252;
wire            n253;
wire            n254;
wire            n255;
wire            n256;
wire            n257;
wire            n258;
wire            n259;
wire            n260;
wire            n261;
wire            n262;
wire            n263;
wire            n264;
wire            n265;
wire      [7:0] n266;
wire      [7:0] n267;
wire      [7:0] n268;
wire      [7:0] n269;
wire      [7:0] n270;
wire      [7:0] n271;
wire      [7:0] n272;
wire      [7:0] n273;
wire      [7:0] n274;
wire      [7:0] n275;
wire            n276;
wire            n277;
wire            n278;
wire            n279;
wire            n280;
wire            n281;
wire            n282;
wire            n283;
wire            n284;
wire            n285;
wire            n286;
wire            n287;
wire            n288;
wire            n289;
wire      [7:0] n290;
wire            n291;
wire      [8:0] n292;
wire      [7:0] n293;
wire            n294;
wire      [7:0] n295;
wire            n296;
wire      [7:0] n297;
wire            n298;
wire      [7:0] n299;
wire            n300;
wire      [7:0] n301;
wire            n302;
wire      [7:0] n303;
wire            n304;
wire      [7:0] n305;
wire      [7:0] n306;
wire      [7:0] n307;
wire      [7:0] n308;
wire      [7:0] n309;
wire      [7:0] n310;
wire      [7:0] n311;
wire      [7:0] n312;
wire      [7:0] n313;
wire      [7:0] n314;
wire      [7:0] n315;
wire      [7:0] n316;
wire      [7:0] n317;
wire      [7:0] n318;
wire      [7:0] n319;
wire      [7:0] n320;
wire      [7:0] n321;
wire      [7:0] n322;
wire      [7:0] n323;
wire      [7:0] n324;
wire      [7:0] n325;
wire      [7:0] n326;
wire      [7:0] n327;
wire      [7:0] n328;
wire      [7:0] n329;
wire      [7:0] n330;
wire      [7:0] n331;
wire      [7:0] n332;
wire      [7:0] n333;
wire      [7:0] n334;
wire      [7:0] n335;
wire      [7:0] n336;
wire      [7:0] n337;
wire      [7:0] n338;
wire      [7:0] n339;
wire      [7:0] n340;
wire      [7:0] n341;
wire      [7:0] n342;
wire      [7:0] n343;
wire      [7:0] n344;
wire      [7:0] n345;
wire      [7:0] n346;
wire      [7:0] n347;
wire      [7:0] n348;
wire      [7:0] n349;
wire      [7:0] n350;
wire      [7:0] n351;
wire      [7:0] n352;
wire      [7:0] n353;
wire      [7:0] n354;
wire      [7:0] n355;
wire      [7:0] n356;
wire      [7:0] n357;
wire      [7:0] n358;
wire      [7:0] n359;
wire      [7:0] n360;
wire      [7:0] n361;
wire      [7:0] n362;
wire     [15:0] n363;
wire     [23:0] n364;
wire     [31:0] n365;
wire     [39:0] n366;
wire     [47:0] n367;
wire     [55:0] n368;
wire     [63:0] n369;
wire     [71:0] n370;
wire     [71:0] n371;
wire     [71:0] n372;
wire     [71:0] n373;
wire     [71:0] n374;
wire     [71:0] n375;
wire     [71:0] n376;
wire     [71:0] n377;
wire     [71:0] n378;
wire     [71:0] n379;
wire     [71:0] n380;
wire     [71:0] n381;
wire     [71:0] n382;
wire            n383;
wire            n384;
wire            n385;
wire            n386;
wire            n387;
wire            n388;
wire            n389;
wire            n390;
wire            n391;
wire            n392;
wire            n393;
wire            n394;
wire            n395;
wire            n396;
wire            n397;
wire            n398;
wire      [7:0] n399;
wire      [7:0] n400;
wire      [7:0] n401;
wire      [7:0] n402;
wire      [7:0] n403;
wire      [7:0] n404;
wire      [7:0] n405;
wire      [7:0] n406;
wire      [7:0] n407;
wire     [15:0] n408;
wire     [23:0] n409;
wire     [31:0] n410;
wire     [39:0] n411;
wire     [47:0] n412;
wire     [55:0] n413;
wire     [63:0] n414;
wire     [71:0] n415;
wire      [7:0] n416;
wire      [7:0] n417;
wire      [7:0] n418;
wire      [7:0] n419;
wire      [7:0] n420;
wire      [7:0] n421;
wire      [7:0] n422;
wire      [7:0] n423;
wire      [7:0] n424;
wire     [15:0] n425;
wire     [23:0] n426;
wire     [31:0] n427;
wire     [39:0] n428;
wire     [47:0] n429;
wire     [55:0] n430;
wire     [63:0] n431;
wire     [71:0] n432;
wire      [7:0] n433;
wire      [7:0] n434;
wire      [7:0] n435;
wire      [7:0] n436;
wire      [7:0] n437;
wire      [7:0] n438;
wire      [7:0] n439;
wire      [7:0] n440;
wire      [7:0] n441;
wire     [15:0] n442;
wire     [23:0] n443;
wire     [31:0] n444;
wire     [39:0] n445;
wire     [47:0] n446;
wire     [55:0] n447;
wire     [63:0] n448;
wire     [71:0] n449;
wire      [7:0] n450;
wire      [7:0] n451;
wire      [7:0] n452;
wire      [7:0] n453;
wire      [7:0] n454;
wire      [7:0] n455;
wire      [7:0] n456;
wire      [7:0] n457;
wire      [7:0] n458;
wire     [15:0] n459;
wire     [23:0] n460;
wire     [31:0] n461;
wire     [39:0] n462;
wire     [47:0] n463;
wire     [55:0] n464;
wire     [63:0] n465;
wire     [71:0] n466;
wire      [7:0] n467;
wire      [7:0] n468;
wire      [7:0] n469;
wire      [7:0] n470;
wire      [7:0] n471;
wire      [7:0] n472;
wire      [7:0] n473;
wire      [7:0] n474;
wire      [7:0] n475;
wire     [15:0] n476;
wire     [23:0] n477;
wire     [31:0] n478;
wire     [39:0] n479;
wire     [47:0] n480;
wire     [55:0] n481;
wire     [63:0] n482;
wire     [71:0] n483;
wire      [7:0] n484;
wire      [7:0] n485;
wire      [7:0] n486;
wire      [7:0] n487;
wire      [7:0] n488;
wire      [7:0] n489;
wire      [7:0] n490;
wire      [7:0] n491;
wire      [7:0] n492;
wire     [15:0] n493;
wire     [23:0] n494;
wire     [31:0] n495;
wire     [39:0] n496;
wire     [47:0] n497;
wire     [55:0] n498;
wire     [63:0] n499;
wire     [71:0] n500;
wire      [7:0] n501;
wire      [7:0] n502;
wire      [7:0] n503;
wire      [7:0] n504;
wire      [7:0] n505;
wire      [7:0] n506;
wire      [7:0] n507;
wire      [7:0] n508;
wire      [7:0] n509;
wire     [15:0] n510;
wire     [23:0] n511;
wire     [31:0] n512;
wire     [39:0] n513;
wire     [47:0] n514;
wire     [55:0] n515;
wire     [63:0] n516;
wire     [71:0] n517;
wire      [7:0] n518;
wire      [7:0] n519;
wire      [7:0] n520;
wire      [7:0] n521;
wire      [7:0] n522;
wire      [7:0] n523;
wire      [7:0] n524;
wire      [7:0] n525;
wire      [7:0] n526;
wire     [15:0] n527;
wire     [23:0] n528;
wire     [31:0] n529;
wire     [39:0] n530;
wire     [47:0] n531;
wire     [55:0] n532;
wire     [63:0] n533;
wire     [71:0] n534;
wire      [7:0] n535;
wire      [7:0] n536;
wire      [7:0] n537;
wire      [7:0] n538;
wire      [7:0] n539;
wire      [7:0] n540;
wire      [7:0] n541;
wire      [7:0] n542;
wire      [7:0] n543;
wire     [15:0] n544;
wire     [23:0] n545;
wire     [31:0] n546;
wire     [39:0] n547;
wire     [47:0] n548;
wire     [55:0] n549;
wire     [63:0] n550;
wire     [71:0] n551;
wire    [143:0] n552;
wire    [215:0] n553;
wire    [287:0] n554;
wire    [359:0] n555;
wire    [431:0] n556;
wire    [503:0] n557;
wire    [575:0] n558;
wire    [647:0] n559;
wire    [647:0] n560;
wire    [647:0] n561;
wire    [647:0] n562;
wire    [647:0] n563;
wire    [647:0] n564;
wire    [647:0] n565;
wire    [647:0] n566;
wire    [647:0] n567;
wire    [647:0] n568;
wire    [647:0] n569;
wire    [647:0] n570;
wire            n571;
wire            n572;
wire            n573;
wire            n574;
wire            n575;
wire            n576;
wire            n577;
wire            n578;
wire            n579;
wire            n580;
wire            n581;
wire            n582;
wire            n583;
wire            n584;
wire            n585;
wire            n586;
wire      [8:0] LB2D_proc_0_addr0;
wire      [7:0] LB2D_proc_0_data0;
wire            n587;
wire            n588;
wire            n589;
wire            n590;
wire            n591;
wire            n592;
wire            n593;
wire            n594;
wire            n595;
wire            n596;
wire            n597;
wire            n598;
wire            n599;
wire            n600;
wire            n601;
wire            n602;
wire      [8:0] LB2D_proc_1_addr0;
wire      [7:0] LB2D_proc_1_data0;
wire            n603;
wire            n604;
wire            n605;
wire      [8:0] LB2D_proc_2_addr0;
wire      [7:0] LB2D_proc_2_data0;
wire            n606;
wire            n607;
wire            n608;
wire      [8:0] LB2D_proc_3_addr0;
wire      [7:0] LB2D_proc_3_data0;
wire            n609;
wire            n610;
wire            n611;
wire      [8:0] LB2D_proc_4_addr0;
wire      [7:0] LB2D_proc_4_data0;
wire            n612;
wire            n613;
wire            n614;
wire      [8:0] LB2D_proc_5_addr0;
wire      [7:0] LB2D_proc_5_data0;
wire            n615;
wire            n616;
wire            n617;
wire      [8:0] LB2D_proc_6_addr0;
wire      [7:0] LB2D_proc_6_data0;
wire            n618;
wire            n619;
wire            n620;
wire      [8:0] LB2D_proc_7_addr0;
wire      [7:0] LB2D_proc_7_data0;
wire            n621;
wire            n622;
wire            n623;
reg      [7:0] LB2D_proc_0[511:0];
reg      [7:0] LB2D_proc_1[511:0];
reg      [7:0] LB2D_proc_2[511:0];
reg      [7:0] LB2D_proc_3[511:0];
reg      [7:0] LB2D_proc_4[511:0];
reg      [7:0] LB2D_proc_5[511:0];
reg      [7:0] LB2D_proc_6[511:0];
reg      [7:0] LB2D_proc_7[511:0];
wire clk;
wire rst;
wire step;
assign n0 =  ( arg_1_TREADY ) == ( 1'd1 )  ;
assign n1 =  ( arg_1_TVALID ) == ( 1'd1 )  ;
assign n2 =  ( n0 ) & ( n1 )  ;
assign n3 =  ( arg_0_TREADY ) == ( 1'd0 )  ;
assign n4 =  ( n2 ) & ( n3 )  ;
assign n5 =  ( arg_0_TVALID ) == ( 1'd0 )  ;
assign n6 =  ( gb_exit_it_1 ) == ( 1'd0 )  ;
assign n7 =  ( stencil_stream_empty ) == ( 1'd0 )  ;
assign n8 =  ( n6 ) & ( n7 )  ;
assign n9 =  ( gb_exit_it_1 ) == ( 1'd1 )  ;
assign n10 =  ( gb_exit_it_8 ) == ( 1'd0 )  ;
assign n11 =  ( n9 ) & ( n10 )  ;
assign n12 =  ( n8 ) | ( n11 )  ;
assign n13 =  ( n5 ) & ( n12 )  ;
assign n14 =  ( slice_stream_empty ) == ( 1'd0 )  ;
assign n15 =  ( LB2D_shift_x ) != ( 9'd488 )  ;
assign n16 =  ( n14 ) & ( n15 )  ;
assign n17 =  ( stencil_stream_full ) == ( 1'd0 )  ;
assign n18 =  ( LB2D_shift_x ) < ( 9'd8 )  ;
assign n19 =  ( n17 ) | ( n18 )  ;
assign n20 =  ( n16 ) & ( n19 )  ;
assign n21 =  ( in_stream_empty ) == ( 1'd0 )  ;
assign n22 =  ( slice_stream_full ) == ( 1'd0 )  ;
assign n23 =  ( LB2D_proc_y ) < ( 10'd8 )  ;
assign n24 =  ( n22 ) | ( n23 )  ;
assign n25 =  ( n21 ) & ( n24 )  ;
assign n26 =  ( arg_1_TREADY ) == ( 1'd0 )  ;
assign n27 =  ( in_stream_full ) == ( 1'd0 )  ;
assign n28 =  ( n26 ) & ( n27 )  ;
assign n29 =  ( LB1D_it_1 ) == ( 1'd0 )  ;
assign n30 =  ( n28 ) & ( n29 )  ;
assign n31 =  ( LB1D_it_1 ) == ( 1'd1 )  ;
assign n32 =  ( n28 ) & ( n31 )  ;
assign n33 =  ( n32 ) ? ( LB1D_uIn ) : ( LB1D_buff ) ;
assign n34 =  ( n30 ) ? ( LB1D_uIn ) : ( n33 ) ;
assign n35 =  ( n25 ) ? ( LB1D_buff ) : ( n34 ) ;
assign n36 =  ( n20 ) ? ( LB1D_buff ) : ( n35 ) ;
assign n37 =  ( n13 ) ? ( LB1D_buff ) : ( n36 ) ;
assign n38 =  ( n4 ) ? ( LB1D_buff ) : ( n37 ) ;
assign n39 =  ( n32 ) ? ( LB1D_in ) : ( LB1D_in ) ;
assign n40 =  ( n30 ) ? ( LB1D_in ) : ( n39 ) ;
assign n41 =  ( n25 ) ? ( LB1D_in ) : ( n40 ) ;
assign n42 =  ( n20 ) ? ( LB1D_in ) : ( n41 ) ;
assign n43 =  ( n13 ) ? ( LB1D_in ) : ( n42 ) ;
assign n44 =  ( n4 ) ? ( arg_1_TDATA ) : ( n43 ) ;
assign n45 =  ( n30 ) ? ( 1'd1 ) : ( LB1D_it_1 ) ;
assign n46 =  ( LB1D_p_cnt ) + ( 19'd1 )  ;
assign n47 =  ( 19'd316224 ) - ( 19'd1 )  ;
assign n48 =  ( LB1D_p_cnt ) == ( n47 )  ;
assign n49 =  ( n48 ) ? ( 19'd0 ) : ( n46 ) ;
assign n50 =  ( n32 ) ? ( n49 ) : ( LB1D_p_cnt ) ;
assign n51 =  ( n30 ) ? ( n46 ) : ( n50 ) ;
assign n52 =  ( n25 ) ? ( LB1D_p_cnt ) : ( n51 ) ;
assign n53 =  ( n20 ) ? ( LB1D_p_cnt ) : ( n52 ) ;
assign n54 =  ( n13 ) ? ( LB1D_p_cnt ) : ( n53 ) ;
assign n55 =  ( n4 ) ? ( LB1D_p_cnt ) : ( n54 ) ;
assign n56 =  ( n32 ) ? ( LB1D_in ) : ( LB1D_uIn ) ;
assign n57 =  ( n30 ) ? ( LB1D_in ) : ( n56 ) ;
assign n58 =  ( n25 ) ? ( LB1D_uIn ) : ( n57 ) ;
assign n59 =  ( n20 ) ? ( LB1D_uIn ) : ( n58 ) ;
assign n60 =  ( n13 ) ? ( LB1D_uIn ) : ( n59 ) ;
assign n61 =  ( n4 ) ? ( LB1D_uIn ) : ( n60 ) ;
assign n62 =  ( LB2D_proc_x ) == ( 9'd488 )  ;
assign n63 =  ( LB2D_proc_w ) == ( 64'd7 )  ;
assign n64 =  ( LB2D_proc_w ) + ( 64'd1 )  ;
assign n65 =  ( n63 ) ? ( 64'd0 ) : ( n64 ) ;
assign n66 =  ( n62 ) ? ( n65 ) : ( LB2D_proc_w ) ;
assign n67 =  ( n32 ) ? ( LB2D_proc_w ) : ( LB2D_proc_w ) ;
assign n68 =  ( n25 ) ? ( n66 ) : ( n67 ) ;
assign n69 =  ( n20 ) ? ( LB2D_proc_w ) : ( n68 ) ;
assign n70 =  ( n13 ) ? ( LB2D_proc_w ) : ( n69 ) ;
assign n71 =  ( n4 ) ? ( LB2D_proc_w ) : ( n70 ) ;
assign n72 =  ( LB2D_proc_x ) + ( 9'd1 )  ;
assign n73 =  ( n62 ) ? ( 9'd1 ) : ( n72 ) ;
assign n74 =  ( n32 ) ? ( LB2D_proc_x ) : ( LB2D_proc_x ) ;
assign n75 =  ( n25 ) ? ( n73 ) : ( n74 ) ;
assign n76 =  ( n20 ) ? ( LB2D_proc_x ) : ( n75 ) ;
assign n77 =  ( n13 ) ? ( LB2D_proc_x ) : ( n76 ) ;
assign n78 =  ( n4 ) ? ( LB2D_proc_x ) : ( n77 ) ;
assign n79 =  ( LB2D_proc_y ) == ( 10'd648 )  ;
assign n80 =  ( LB2D_proc_y ) + ( 10'd1 )  ;
assign n81 =  ( n79 ) ? ( 10'd0 ) : ( n80 ) ;
assign n82 =  ( n62 ) ? ( n81 ) : ( LB2D_proc_y ) ;
assign n83 =  ( n32 ) ? ( LB2D_proc_y ) : ( LB2D_proc_y ) ;
assign n84 =  ( n25 ) ? ( n82 ) : ( n83 ) ;
assign n85 =  ( n20 ) ? ( LB2D_proc_y ) : ( n84 ) ;
assign n86 =  ( n13 ) ? ( LB2D_proc_y ) : ( n85 ) ;
assign n87 =  ( n4 ) ? ( LB2D_proc_y ) : ( n86 ) ;
assign n88 =  ( n32 ) ? ( LB2D_shift_0 ) : ( LB2D_shift_0 ) ;
assign n89 =  ( n25 ) ? ( LB2D_shift_0 ) : ( n88 ) ;
assign n90 =  ( n20 ) ? ( LB2D_shift_1 ) : ( n89 ) ;
assign n91 =  ( n13 ) ? ( LB2D_shift_0 ) : ( n90 ) ;
assign n92 =  ( n4 ) ? ( LB2D_shift_0 ) : ( n91 ) ;
assign n93 =  ( n32 ) ? ( LB2D_shift_1 ) : ( LB2D_shift_1 ) ;
assign n94 =  ( n25 ) ? ( LB2D_shift_1 ) : ( n93 ) ;
assign n95 =  ( n20 ) ? ( LB2D_shift_2 ) : ( n94 ) ;
assign n96 =  ( n13 ) ? ( LB2D_shift_1 ) : ( n95 ) ;
assign n97 =  ( n4 ) ? ( LB2D_shift_1 ) : ( n96 ) ;
assign n98 =  ( n32 ) ? ( LB2D_shift_2 ) : ( LB2D_shift_2 ) ;
assign n99 =  ( n25 ) ? ( LB2D_shift_2 ) : ( n98 ) ;
assign n100 =  ( n20 ) ? ( LB2D_shift_3 ) : ( n99 ) ;
assign n101 =  ( n13 ) ? ( LB2D_shift_2 ) : ( n100 ) ;
assign n102 =  ( n4 ) ? ( LB2D_shift_2 ) : ( n101 ) ;
assign n103 =  ( n32 ) ? ( LB2D_shift_3 ) : ( LB2D_shift_3 ) ;
assign n104 =  ( n25 ) ? ( LB2D_shift_3 ) : ( n103 ) ;
assign n105 =  ( n20 ) ? ( LB2D_shift_4 ) : ( n104 ) ;
assign n106 =  ( n13 ) ? ( LB2D_shift_3 ) : ( n105 ) ;
assign n107 =  ( n4 ) ? ( LB2D_shift_3 ) : ( n106 ) ;
assign n108 =  ( n32 ) ? ( LB2D_shift_4 ) : ( LB2D_shift_4 ) ;
assign n109 =  ( n25 ) ? ( LB2D_shift_4 ) : ( n108 ) ;
assign n110 =  ( n20 ) ? ( LB2D_shift_5 ) : ( n109 ) ;
assign n111 =  ( n13 ) ? ( LB2D_shift_4 ) : ( n110 ) ;
assign n112 =  ( n4 ) ? ( LB2D_shift_4 ) : ( n111 ) ;
assign n113 =  ( n32 ) ? ( LB2D_shift_5 ) : ( LB2D_shift_5 ) ;
assign n114 =  ( n25 ) ? ( LB2D_shift_5 ) : ( n113 ) ;
assign n115 =  ( n20 ) ? ( LB2D_shift_6 ) : ( n114 ) ;
assign n116 =  ( n13 ) ? ( LB2D_shift_5 ) : ( n115 ) ;
assign n117 =  ( n4 ) ? ( LB2D_shift_5 ) : ( n116 ) ;
assign n118 =  ( n32 ) ? ( LB2D_shift_6 ) : ( LB2D_shift_6 ) ;
assign n119 =  ( n25 ) ? ( LB2D_shift_6 ) : ( n118 ) ;
assign n120 =  ( n20 ) ? ( LB2D_shift_7 ) : ( n119 ) ;
assign n121 =  ( n13 ) ? ( LB2D_shift_6 ) : ( n120 ) ;
assign n122 =  ( n4 ) ? ( LB2D_shift_6 ) : ( n121 ) ;
assign n123 =  ( slice_stream_full ) == ( 1'd1 )  ;
assign n124 =  ( n123 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n125 =  ( n32 ) ? ( LB2D_shift_7 ) : ( LB2D_shift_7 ) ;
assign n126 =  ( n25 ) ? ( LB2D_shift_7 ) : ( n125 ) ;
assign n127 =  ( n20 ) ? ( n124 ) : ( n126 ) ;
assign n128 =  ( n13 ) ? ( LB2D_shift_7 ) : ( n127 ) ;
assign n129 =  ( n4 ) ? ( LB2D_shift_7 ) : ( n128 ) ;
assign n130 =  ( LB2D_shift_x ) == ( 9'd488 )  ;
assign n131 =  ( n14 ) & ( n130 )  ;
assign n132 =  ( n131 ) & ( n19 )  ;
assign n133 =  ( LB2D_shift_x ) + ( 9'd1 )  ;
assign n134 =  ( n32 ) ? ( LB2D_shift_x ) : ( LB2D_shift_x ) ;
assign n135 =  ( n25 ) ? ( LB2D_shift_x ) : ( n134 ) ;
assign n136 =  ( n20 ) ? ( n133 ) : ( n135 ) ;
assign n137 =  ( n132 ) ? ( 9'd0 ) : ( n136 ) ;
assign n138 =  ( n13 ) ? ( LB2D_shift_x ) : ( n137 ) ;
assign n139 =  ( n4 ) ? ( LB2D_shift_x ) : ( n138 ) ;
assign n140 =  ( LB2D_shift_y ) < ( 10'd640 )  ;
assign n141 =  ( LB2D_shift_x ) < ( 9'd488 )  ;
assign n142 =  ( LB2D_shift_y ) + ( 10'd1 )  ;
assign n143 =  ( n141 ) ? ( LB2D_shift_y ) : ( n142 ) ;
assign n144 =  ( n140 ) ? ( n143 ) : ( 10'd640 ) ;
assign n145 =  ( n32 ) ? ( LB2D_shift_y ) : ( LB2D_shift_y ) ;
assign n146 =  ( n25 ) ? ( LB2D_shift_y ) : ( n145 ) ;
assign n147 =  ( n20 ) ? ( n144 ) : ( n146 ) ;
assign n148 =  ( n13 ) ? ( LB2D_shift_y ) : ( n147 ) ;
assign n149 =  ( n4 ) ? ( LB2D_shift_y ) : ( n148 ) ;
assign n150 =  ( stencil_stream_full ) == ( 1'd1 )  ;
assign n151 =  ( n150 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_0 ) ;
assign n152 = gb_fun(n151) ;
assign n153 =  ( n32 ) ? ( arg_0_TDATA ) : ( arg_0_TDATA ) ;
assign n154 =  ( n25 ) ? ( arg_0_TDATA ) : ( n153 ) ;
assign n155 =  ( n20 ) ? ( arg_0_TDATA ) : ( n154 ) ;
assign n156 =  ( n13 ) ? ( n152 ) : ( n155 ) ;
assign n157 =  ( n4 ) ? ( arg_0_TDATA ) : ( n156 ) ;
assign n158 =  ( gb_pp_it_8 ) == ( 1'd1 )  ;
assign n159 =  ( n158 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n160 =  ( n32 ) ? ( arg_0_TVALID ) : ( arg_0_TVALID ) ;
assign n161 =  ( n25 ) ? ( arg_0_TVALID ) : ( n160 ) ;
assign n162 =  ( n20 ) ? ( arg_0_TVALID ) : ( n161 ) ;
assign n163 =  ( n13 ) ? ( n159 ) : ( n162 ) ;
assign n164 =  ( n4 ) ? ( arg_0_TVALID ) : ( n163 ) ;
assign n165 =  ( n32 ) ? ( 1'd1 ) : ( arg_1_TREADY ) ;
assign n166 =  ( n30 ) ? ( 1'd1 ) : ( n165 ) ;
assign n167 =  ( n25 ) ? ( arg_1_TREADY ) : ( n166 ) ;
assign n168 =  ( n20 ) ? ( arg_1_TREADY ) : ( n167 ) ;
assign n169 =  ( n13 ) ? ( arg_1_TREADY ) : ( n168 ) ;
assign n170 =  ( n4 ) ? ( 1'd0 ) : ( n169 ) ;
assign n171 =  ( gb_p_cnt ) + ( 19'd1 )  ;
assign n172 =  ( n171 ) == ( 19'd307200 )  ;
assign n173 =  ( n172 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n174 =  ( n32 ) ? ( gb_exit_it_1 ) : ( gb_exit_it_1 ) ;
assign n175 =  ( n25 ) ? ( gb_exit_it_1 ) : ( n174 ) ;
assign n176 =  ( n20 ) ? ( gb_exit_it_1 ) : ( n175 ) ;
assign n177 =  ( n13 ) ? ( n173 ) : ( n176 ) ;
assign n178 =  ( n4 ) ? ( gb_exit_it_1 ) : ( n177 ) ;
assign n179 =  ( n32 ) ? ( gb_exit_it_2 ) : ( gb_exit_it_2 ) ;
assign n180 =  ( n25 ) ? ( gb_exit_it_2 ) : ( n179 ) ;
assign n181 =  ( n20 ) ? ( gb_exit_it_2 ) : ( n180 ) ;
assign n182 =  ( n13 ) ? ( gb_exit_it_1 ) : ( n181 ) ;
assign n183 =  ( n4 ) ? ( gb_exit_it_2 ) : ( n182 ) ;
assign n184 =  ( n32 ) ? ( gb_exit_it_3 ) : ( gb_exit_it_3 ) ;
assign n185 =  ( n25 ) ? ( gb_exit_it_3 ) : ( n184 ) ;
assign n186 =  ( n20 ) ? ( gb_exit_it_3 ) : ( n185 ) ;
assign n187 =  ( n13 ) ? ( gb_exit_it_2 ) : ( n186 ) ;
assign n188 =  ( n4 ) ? ( gb_exit_it_3 ) : ( n187 ) ;
assign n189 =  ( n32 ) ? ( gb_exit_it_4 ) : ( gb_exit_it_4 ) ;
assign n190 =  ( n25 ) ? ( gb_exit_it_4 ) : ( n189 ) ;
assign n191 =  ( n20 ) ? ( gb_exit_it_4 ) : ( n190 ) ;
assign n192 =  ( n13 ) ? ( gb_exit_it_3 ) : ( n191 ) ;
assign n193 =  ( n4 ) ? ( gb_exit_it_4 ) : ( n192 ) ;
assign n194 =  ( n32 ) ? ( gb_exit_it_5 ) : ( gb_exit_it_5 ) ;
assign n195 =  ( n25 ) ? ( gb_exit_it_5 ) : ( n194 ) ;
assign n196 =  ( n20 ) ? ( gb_exit_it_5 ) : ( n195 ) ;
assign n197 =  ( n13 ) ? ( gb_exit_it_4 ) : ( n196 ) ;
assign n198 =  ( n4 ) ? ( gb_exit_it_5 ) : ( n197 ) ;
assign n199 =  ( n32 ) ? ( gb_exit_it_6 ) : ( gb_exit_it_6 ) ;
assign n200 =  ( n25 ) ? ( gb_exit_it_6 ) : ( n199 ) ;
assign n201 =  ( n20 ) ? ( gb_exit_it_6 ) : ( n200 ) ;
assign n202 =  ( n13 ) ? ( gb_exit_it_5 ) : ( n201 ) ;
assign n203 =  ( n4 ) ? ( gb_exit_it_6 ) : ( n202 ) ;
assign n204 =  ( n32 ) ? ( gb_exit_it_7 ) : ( gb_exit_it_7 ) ;
assign n205 =  ( n25 ) ? ( gb_exit_it_7 ) : ( n204 ) ;
assign n206 =  ( n20 ) ? ( gb_exit_it_7 ) : ( n205 ) ;
assign n207 =  ( n13 ) ? ( gb_exit_it_6 ) : ( n206 ) ;
assign n208 =  ( n4 ) ? ( gb_exit_it_7 ) : ( n207 ) ;
assign n209 =  ( n32 ) ? ( gb_exit_it_8 ) : ( gb_exit_it_8 ) ;
assign n210 =  ( n25 ) ? ( gb_exit_it_8 ) : ( n209 ) ;
assign n211 =  ( n20 ) ? ( gb_exit_it_8 ) : ( n210 ) ;
assign n212 =  ( n13 ) ? ( gb_exit_it_7 ) : ( n211 ) ;
assign n213 =  ( n4 ) ? ( gb_exit_it_8 ) : ( n212 ) ;
assign n214 =  ( gb_p_cnt ) < ( 19'd307200 )  ;
assign n215 =  ( n214 ) ? ( n171 ) : ( 19'd307200 ) ;
assign n216 =  ( n32 ) ? ( gb_p_cnt ) : ( gb_p_cnt ) ;
assign n217 =  ( n25 ) ? ( gb_p_cnt ) : ( n216 ) ;
assign n218 =  ( n20 ) ? ( gb_p_cnt ) : ( n217 ) ;
assign n219 =  ( n13 ) ? ( n215 ) : ( n218 ) ;
assign n220 =  ( n4 ) ? ( gb_p_cnt ) : ( n219 ) ;
assign n221 =  ( n32 ) ? ( gb_pp_it_1 ) : ( gb_pp_it_1 ) ;
assign n222 =  ( n25 ) ? ( gb_pp_it_1 ) : ( n221 ) ;
assign n223 =  ( n20 ) ? ( gb_pp_it_1 ) : ( n222 ) ;
assign n224 =  ( n13 ) ? ( 1'd1 ) : ( n223 ) ;
assign n225 =  ( n4 ) ? ( gb_pp_it_1 ) : ( n224 ) ;
assign n226 =  ( n32 ) ? ( gb_pp_it_2 ) : ( gb_pp_it_2 ) ;
assign n227 =  ( n25 ) ? ( gb_pp_it_2 ) : ( n226 ) ;
assign n228 =  ( n20 ) ? ( gb_pp_it_2 ) : ( n227 ) ;
assign n229 =  ( n13 ) ? ( gb_pp_it_1 ) : ( n228 ) ;
assign n230 =  ( n4 ) ? ( gb_pp_it_2 ) : ( n229 ) ;
assign n231 =  ( n32 ) ? ( gb_pp_it_3 ) : ( gb_pp_it_3 ) ;
assign n232 =  ( n25 ) ? ( gb_pp_it_3 ) : ( n231 ) ;
assign n233 =  ( n20 ) ? ( gb_pp_it_3 ) : ( n232 ) ;
assign n234 =  ( n13 ) ? ( gb_pp_it_2 ) : ( n233 ) ;
assign n235 =  ( n4 ) ? ( gb_pp_it_3 ) : ( n234 ) ;
assign n236 =  ( n32 ) ? ( gb_pp_it_4 ) : ( gb_pp_it_4 ) ;
assign n237 =  ( n25 ) ? ( gb_pp_it_4 ) : ( n236 ) ;
assign n238 =  ( n20 ) ? ( gb_pp_it_4 ) : ( n237 ) ;
assign n239 =  ( n13 ) ? ( gb_pp_it_3 ) : ( n238 ) ;
assign n240 =  ( n4 ) ? ( gb_pp_it_4 ) : ( n239 ) ;
assign n241 =  ( n32 ) ? ( gb_pp_it_5 ) : ( gb_pp_it_5 ) ;
assign n242 =  ( n25 ) ? ( gb_pp_it_5 ) : ( n241 ) ;
assign n243 =  ( n20 ) ? ( gb_pp_it_5 ) : ( n242 ) ;
assign n244 =  ( n13 ) ? ( gb_pp_it_4 ) : ( n243 ) ;
assign n245 =  ( n4 ) ? ( gb_pp_it_5 ) : ( n244 ) ;
assign n246 =  ( n32 ) ? ( gb_pp_it_6 ) : ( gb_pp_it_6 ) ;
assign n247 =  ( n25 ) ? ( gb_pp_it_6 ) : ( n246 ) ;
assign n248 =  ( n20 ) ? ( gb_pp_it_6 ) : ( n247 ) ;
assign n249 =  ( n13 ) ? ( gb_pp_it_5 ) : ( n248 ) ;
assign n250 =  ( n4 ) ? ( gb_pp_it_6 ) : ( n249 ) ;
assign n251 =  ( n32 ) ? ( gb_pp_it_7 ) : ( gb_pp_it_7 ) ;
assign n252 =  ( n25 ) ? ( gb_pp_it_7 ) : ( n251 ) ;
assign n253 =  ( n20 ) ? ( gb_pp_it_7 ) : ( n252 ) ;
assign n254 =  ( n13 ) ? ( gb_pp_it_6 ) : ( n253 ) ;
assign n255 =  ( n4 ) ? ( gb_pp_it_7 ) : ( n254 ) ;
assign n256 =  ( n32 ) ? ( gb_pp_it_8 ) : ( gb_pp_it_8 ) ;
assign n257 =  ( n25 ) ? ( gb_pp_it_8 ) : ( n256 ) ;
assign n258 =  ( n20 ) ? ( gb_pp_it_8 ) : ( n257 ) ;
assign n259 =  ( n13 ) ? ( gb_pp_it_7 ) : ( n258 ) ;
assign n260 =  ( n4 ) ? ( gb_pp_it_8 ) : ( n259 ) ;
assign n261 =  ( n32 ) ? ( gb_pp_it_9 ) : ( gb_pp_it_9 ) ;
assign n262 =  ( n25 ) ? ( gb_pp_it_9 ) : ( n261 ) ;
assign n263 =  ( n20 ) ? ( gb_pp_it_9 ) : ( n262 ) ;
assign n264 =  ( n13 ) ? ( gb_pp_it_8 ) : ( n263 ) ;
assign n265 =  ( n4 ) ? ( gb_pp_it_9 ) : ( n264 ) ;
assign n266 =  ( n32 ) ? ( LB1D_buff ) : ( in_stream_buff_0 ) ;
assign n267 =  ( n25 ) ? ( in_stream_buff_0 ) : ( n266 ) ;
assign n268 =  ( n20 ) ? ( in_stream_buff_0 ) : ( n267 ) ;
assign n269 =  ( n13 ) ? ( in_stream_buff_0 ) : ( n268 ) ;
assign n270 =  ( n4 ) ? ( in_stream_buff_0 ) : ( n269 ) ;
assign n271 =  ( n32 ) ? ( in_stream_buff_0 ) : ( in_stream_buff_1 ) ;
assign n272 =  ( n25 ) ? ( in_stream_buff_1 ) : ( n271 ) ;
assign n273 =  ( n20 ) ? ( in_stream_buff_1 ) : ( n272 ) ;
assign n274 =  ( n13 ) ? ( in_stream_buff_1 ) : ( n273 ) ;
assign n275 =  ( n4 ) ? ( in_stream_buff_1 ) : ( n274 ) ;
assign n276 =  ( in_stream_full ) == ( 1'd1 )  ;
assign n277 =  ( n276 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n278 =  ( n32 ) ? ( 1'd0 ) : ( in_stream_empty ) ;
assign n279 =  ( n25 ) ? ( n277 ) : ( n278 ) ;
assign n280 =  ( n20 ) ? ( in_stream_empty ) : ( n279 ) ;
assign n281 =  ( n13 ) ? ( in_stream_empty ) : ( n280 ) ;
assign n282 =  ( n4 ) ? ( in_stream_empty ) : ( n281 ) ;
assign n283 =  ( in_stream_empty ) == ( 1'd1 )  ;
assign n284 =  ( n283 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n285 =  ( n32 ) ? ( n284 ) : ( in_stream_full ) ;
assign n286 =  ( n25 ) ? ( 1'd0 ) : ( n285 ) ;
assign n287 =  ( n20 ) ? ( in_stream_full ) : ( n286 ) ;
assign n288 =  ( n13 ) ? ( in_stream_full ) : ( n287 ) ;
assign n289 =  ( n4 ) ? ( in_stream_full ) : ( n288 ) ;
assign n290 =  ( n276 ) ? ( in_stream_buff_1 ) : ( in_stream_buff_0 ) ;
assign n291 =  ( LB2D_proc_w ) == ( 64'd0 )  ;
assign n292 =  ( LB2D_proc_x ) - ( 9'd1 )  ;
assign n293 =  (  LB2D_proc_7 [ n292 ] )  ;
assign n294 =  ( LB2D_proc_w ) == ( 64'd1 )  ;
assign n295 =  (  LB2D_proc_0 [ n292 ] )  ;
assign n296 =  ( LB2D_proc_w ) == ( 64'd2 )  ;
assign n297 =  (  LB2D_proc_1 [ n292 ] )  ;
assign n298 =  ( LB2D_proc_w ) == ( 64'd3 )  ;
assign n299 =  (  LB2D_proc_2 [ n292 ] )  ;
assign n300 =  ( LB2D_proc_w ) == ( 64'd4 )  ;
assign n301 =  (  LB2D_proc_3 [ n292 ] )  ;
assign n302 =  ( LB2D_proc_w ) == ( 64'd5 )  ;
assign n303 =  (  LB2D_proc_4 [ n292 ] )  ;
assign n304 =  ( LB2D_proc_w ) == ( 64'd6 )  ;
assign n305 =  (  LB2D_proc_5 [ n292 ] )  ;
assign n306 =  (  LB2D_proc_6 [ n292 ] )  ;
assign n307 =  ( n304 ) ? ( n305 ) : ( n306 ) ;
assign n308 =  ( n302 ) ? ( n303 ) : ( n307 ) ;
assign n309 =  ( n300 ) ? ( n301 ) : ( n308 ) ;
assign n310 =  ( n298 ) ? ( n299 ) : ( n309 ) ;
assign n311 =  ( n296 ) ? ( n297 ) : ( n310 ) ;
assign n312 =  ( n294 ) ? ( n295 ) : ( n311 ) ;
assign n313 =  ( n291 ) ? ( n293 ) : ( n312 ) ;
assign n314 =  ( n304 ) ? ( n303 ) : ( n305 ) ;
assign n315 =  ( n302 ) ? ( n301 ) : ( n314 ) ;
assign n316 =  ( n300 ) ? ( n299 ) : ( n315 ) ;
assign n317 =  ( n298 ) ? ( n297 ) : ( n316 ) ;
assign n318 =  ( n296 ) ? ( n295 ) : ( n317 ) ;
assign n319 =  ( n294 ) ? ( n293 ) : ( n318 ) ;
assign n320 =  ( n291 ) ? ( n306 ) : ( n319 ) ;
assign n321 =  ( n304 ) ? ( n301 ) : ( n303 ) ;
assign n322 =  ( n302 ) ? ( n299 ) : ( n321 ) ;
assign n323 =  ( n300 ) ? ( n297 ) : ( n322 ) ;
assign n324 =  ( n298 ) ? ( n295 ) : ( n323 ) ;
assign n325 =  ( n296 ) ? ( n293 ) : ( n324 ) ;
assign n326 =  ( n294 ) ? ( n306 ) : ( n325 ) ;
assign n327 =  ( n291 ) ? ( n305 ) : ( n326 ) ;
assign n328 =  ( n304 ) ? ( n299 ) : ( n301 ) ;
assign n329 =  ( n302 ) ? ( n297 ) : ( n328 ) ;
assign n330 =  ( n300 ) ? ( n295 ) : ( n329 ) ;
assign n331 =  ( n298 ) ? ( n293 ) : ( n330 ) ;
assign n332 =  ( n296 ) ? ( n306 ) : ( n331 ) ;
assign n333 =  ( n294 ) ? ( n305 ) : ( n332 ) ;
assign n334 =  ( n291 ) ? ( n303 ) : ( n333 ) ;
assign n335 =  ( n304 ) ? ( n297 ) : ( n299 ) ;
assign n336 =  ( n302 ) ? ( n295 ) : ( n335 ) ;
assign n337 =  ( n300 ) ? ( n293 ) : ( n336 ) ;
assign n338 =  ( n298 ) ? ( n306 ) : ( n337 ) ;
assign n339 =  ( n296 ) ? ( n305 ) : ( n338 ) ;
assign n340 =  ( n294 ) ? ( n303 ) : ( n339 ) ;
assign n341 =  ( n291 ) ? ( n301 ) : ( n340 ) ;
assign n342 =  ( n304 ) ? ( n295 ) : ( n297 ) ;
assign n343 =  ( n302 ) ? ( n293 ) : ( n342 ) ;
assign n344 =  ( n300 ) ? ( n306 ) : ( n343 ) ;
assign n345 =  ( n298 ) ? ( n305 ) : ( n344 ) ;
assign n346 =  ( n296 ) ? ( n303 ) : ( n345 ) ;
assign n347 =  ( n294 ) ? ( n301 ) : ( n346 ) ;
assign n348 =  ( n291 ) ? ( n299 ) : ( n347 ) ;
assign n349 =  ( n304 ) ? ( n293 ) : ( n295 ) ;
assign n350 =  ( n302 ) ? ( n306 ) : ( n349 ) ;
assign n351 =  ( n300 ) ? ( n305 ) : ( n350 ) ;
assign n352 =  ( n298 ) ? ( n303 ) : ( n351 ) ;
assign n353 =  ( n296 ) ? ( n301 ) : ( n352 ) ;
assign n354 =  ( n294 ) ? ( n299 ) : ( n353 ) ;
assign n355 =  ( n291 ) ? ( n297 ) : ( n354 ) ;
assign n356 =  ( n304 ) ? ( n306 ) : ( n293 ) ;
assign n357 =  ( n302 ) ? ( n305 ) : ( n356 ) ;
assign n358 =  ( n300 ) ? ( n303 ) : ( n357 ) ;
assign n359 =  ( n298 ) ? ( n301 ) : ( n358 ) ;
assign n360 =  ( n296 ) ? ( n299 ) : ( n359 ) ;
assign n361 =  ( n294 ) ? ( n297 ) : ( n360 ) ;
assign n362 =  ( n291 ) ? ( n295 ) : ( n361 ) ;
assign n363 =  { ( n355 ) , ( n362 ) }  ;
assign n364 =  { ( n348 ) , ( n363 ) }  ;
assign n365 =  { ( n341 ) , ( n364 ) }  ;
assign n366 =  { ( n334 ) , ( n365 ) }  ;
assign n367 =  { ( n327 ) , ( n366 ) }  ;
assign n368 =  { ( n320 ) , ( n367 ) }  ;
assign n369 =  { ( n313 ) , ( n368 ) }  ;
assign n370 =  { ( n290 ) , ( n369 ) }  ;
assign n371 =  ( n23 ) ? ( slice_stream_buff_0 ) : ( n370 ) ;
assign n372 =  ( n32 ) ? ( slice_stream_buff_0 ) : ( slice_stream_buff_0 ) ;
assign n373 =  ( n25 ) ? ( n371 ) : ( n372 ) ;
assign n374 =  ( n20 ) ? ( slice_stream_buff_0 ) : ( n373 ) ;
assign n375 =  ( n13 ) ? ( slice_stream_buff_0 ) : ( n374 ) ;
assign n376 =  ( n4 ) ? ( slice_stream_buff_0 ) : ( n375 ) ;
assign n377 =  ( n23 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n378 =  ( n32 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_1 ) ;
assign n379 =  ( n25 ) ? ( n377 ) : ( n378 ) ;
assign n380 =  ( n20 ) ? ( slice_stream_buff_1 ) : ( n379 ) ;
assign n381 =  ( n13 ) ? ( slice_stream_buff_1 ) : ( n380 ) ;
assign n382 =  ( n4 ) ? ( slice_stream_buff_1 ) : ( n381 ) ;
assign n383 =  ( n123 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n384 =  ( n23 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n385 =  ( n32 ) ? ( slice_stream_empty ) : ( slice_stream_empty ) ;
assign n386 =  ( n25 ) ? ( n384 ) : ( n385 ) ;
assign n387 =  ( n20 ) ? ( n383 ) : ( n386 ) ;
assign n388 =  ( n13 ) ? ( slice_stream_empty ) : ( n387 ) ;
assign n389 =  ( n4 ) ? ( slice_stream_empty ) : ( n388 ) ;
assign n390 =  ( slice_stream_empty ) == ( 1'd1 )  ;
assign n391 =  ( n390 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n392 =  ( n23 ) ? ( 1'd0 ) : ( n391 ) ;
assign n393 =  ( n32 ) ? ( slice_stream_full ) : ( slice_stream_full ) ;
assign n394 =  ( n25 ) ? ( n392 ) : ( n393 ) ;
assign n395 =  ( n20 ) ? ( 1'd0 ) : ( n394 ) ;
assign n396 =  ( n13 ) ? ( slice_stream_full ) : ( n395 ) ;
assign n397 =  ( n4 ) ? ( slice_stream_full ) : ( n396 ) ;
assign n398 =  ( LB2D_shift_x ) >= ( 9'd8 )  ;
assign n399 = n124[71:64] ;
assign n400 = LB2D_shift_7[71:64] ;
assign n401 = LB2D_shift_6[71:64] ;
assign n402 = LB2D_shift_5[71:64] ;
assign n403 = LB2D_shift_4[71:64] ;
assign n404 = LB2D_shift_3[71:64] ;
assign n405 = LB2D_shift_2[71:64] ;
assign n406 = LB2D_shift_1[71:64] ;
assign n407 = LB2D_shift_0[71:64] ;
assign n408 =  { ( n406 ) , ( n407 ) }  ;
assign n409 =  { ( n405 ) , ( n408 ) }  ;
assign n410 =  { ( n404 ) , ( n409 ) }  ;
assign n411 =  { ( n403 ) , ( n410 ) }  ;
assign n412 =  { ( n402 ) , ( n411 ) }  ;
assign n413 =  { ( n401 ) , ( n412 ) }  ;
assign n414 =  { ( n400 ) , ( n413 ) }  ;
assign n415 =  { ( n399 ) , ( n414 ) }  ;
assign n416 = n124[63:56] ;
assign n417 = LB2D_shift_7[63:56] ;
assign n418 = LB2D_shift_6[63:56] ;
assign n419 = LB2D_shift_5[63:56] ;
assign n420 = LB2D_shift_4[63:56] ;
assign n421 = LB2D_shift_3[63:56] ;
assign n422 = LB2D_shift_2[63:56] ;
assign n423 = LB2D_shift_1[63:56] ;
assign n424 = LB2D_shift_0[63:56] ;
assign n425 =  { ( n423 ) , ( n424 ) }  ;
assign n426 =  { ( n422 ) , ( n425 ) }  ;
assign n427 =  { ( n421 ) , ( n426 ) }  ;
assign n428 =  { ( n420 ) , ( n427 ) }  ;
assign n429 =  { ( n419 ) , ( n428 ) }  ;
assign n430 =  { ( n418 ) , ( n429 ) }  ;
assign n431 =  { ( n417 ) , ( n430 ) }  ;
assign n432 =  { ( n416 ) , ( n431 ) }  ;
assign n433 = n124[55:48] ;
assign n434 = LB2D_shift_7[55:48] ;
assign n435 = LB2D_shift_6[55:48] ;
assign n436 = LB2D_shift_5[55:48] ;
assign n437 = LB2D_shift_4[55:48] ;
assign n438 = LB2D_shift_3[55:48] ;
assign n439 = LB2D_shift_2[55:48] ;
assign n440 = LB2D_shift_1[55:48] ;
assign n441 = LB2D_shift_0[55:48] ;
assign n442 =  { ( n440 ) , ( n441 ) }  ;
assign n443 =  { ( n439 ) , ( n442 ) }  ;
assign n444 =  { ( n438 ) , ( n443 ) }  ;
assign n445 =  { ( n437 ) , ( n444 ) }  ;
assign n446 =  { ( n436 ) , ( n445 ) }  ;
assign n447 =  { ( n435 ) , ( n446 ) }  ;
assign n448 =  { ( n434 ) , ( n447 ) }  ;
assign n449 =  { ( n433 ) , ( n448 ) }  ;
assign n450 = n124[47:40] ;
assign n451 = LB2D_shift_7[47:40] ;
assign n452 = LB2D_shift_6[47:40] ;
assign n453 = LB2D_shift_5[47:40] ;
assign n454 = LB2D_shift_4[47:40] ;
assign n455 = LB2D_shift_3[47:40] ;
assign n456 = LB2D_shift_2[47:40] ;
assign n457 = LB2D_shift_1[47:40] ;
assign n458 = LB2D_shift_0[47:40] ;
assign n459 =  { ( n457 ) , ( n458 ) }  ;
assign n460 =  { ( n456 ) , ( n459 ) }  ;
assign n461 =  { ( n455 ) , ( n460 ) }  ;
assign n462 =  { ( n454 ) , ( n461 ) }  ;
assign n463 =  { ( n453 ) , ( n462 ) }  ;
assign n464 =  { ( n452 ) , ( n463 ) }  ;
assign n465 =  { ( n451 ) , ( n464 ) }  ;
assign n466 =  { ( n450 ) , ( n465 ) }  ;
assign n467 = n124[39:32] ;
assign n468 = LB2D_shift_7[39:32] ;
assign n469 = LB2D_shift_6[39:32] ;
assign n470 = LB2D_shift_5[39:32] ;
assign n471 = LB2D_shift_4[39:32] ;
assign n472 = LB2D_shift_3[39:32] ;
assign n473 = LB2D_shift_2[39:32] ;
assign n474 = LB2D_shift_1[39:32] ;
assign n475 = LB2D_shift_0[39:32] ;
assign n476 =  { ( n474 ) , ( n475 ) }  ;
assign n477 =  { ( n473 ) , ( n476 ) }  ;
assign n478 =  { ( n472 ) , ( n477 ) }  ;
assign n479 =  { ( n471 ) , ( n478 ) }  ;
assign n480 =  { ( n470 ) , ( n479 ) }  ;
assign n481 =  { ( n469 ) , ( n480 ) }  ;
assign n482 =  { ( n468 ) , ( n481 ) }  ;
assign n483 =  { ( n467 ) , ( n482 ) }  ;
assign n484 = n124[31:24] ;
assign n485 = LB2D_shift_7[31:24] ;
assign n486 = LB2D_shift_6[31:24] ;
assign n487 = LB2D_shift_5[31:24] ;
assign n488 = LB2D_shift_4[31:24] ;
assign n489 = LB2D_shift_3[31:24] ;
assign n490 = LB2D_shift_2[31:24] ;
assign n491 = LB2D_shift_1[31:24] ;
assign n492 = LB2D_shift_0[31:24] ;
assign n493 =  { ( n491 ) , ( n492 ) }  ;
assign n494 =  { ( n490 ) , ( n493 ) }  ;
assign n495 =  { ( n489 ) , ( n494 ) }  ;
assign n496 =  { ( n488 ) , ( n495 ) }  ;
assign n497 =  { ( n487 ) , ( n496 ) }  ;
assign n498 =  { ( n486 ) , ( n497 ) }  ;
assign n499 =  { ( n485 ) , ( n498 ) }  ;
assign n500 =  { ( n484 ) , ( n499 ) }  ;
assign n501 = n124[23:16] ;
assign n502 = LB2D_shift_7[23:16] ;
assign n503 = LB2D_shift_6[23:16] ;
assign n504 = LB2D_shift_5[23:16] ;
assign n505 = LB2D_shift_4[23:16] ;
assign n506 = LB2D_shift_3[23:16] ;
assign n507 = LB2D_shift_2[23:16] ;
assign n508 = LB2D_shift_1[23:16] ;
assign n509 = LB2D_shift_0[23:16] ;
assign n510 =  { ( n508 ) , ( n509 ) }  ;
assign n511 =  { ( n507 ) , ( n510 ) }  ;
assign n512 =  { ( n506 ) , ( n511 ) }  ;
assign n513 =  { ( n505 ) , ( n512 ) }  ;
assign n514 =  { ( n504 ) , ( n513 ) }  ;
assign n515 =  { ( n503 ) , ( n514 ) }  ;
assign n516 =  { ( n502 ) , ( n515 ) }  ;
assign n517 =  { ( n501 ) , ( n516 ) }  ;
assign n518 = n124[15:8] ;
assign n519 = LB2D_shift_7[15:8] ;
assign n520 = LB2D_shift_6[15:8] ;
assign n521 = LB2D_shift_5[15:8] ;
assign n522 = LB2D_shift_4[15:8] ;
assign n523 = LB2D_shift_3[15:8] ;
assign n524 = LB2D_shift_2[15:8] ;
assign n525 = LB2D_shift_1[15:8] ;
assign n526 = LB2D_shift_0[15:8] ;
assign n527 =  { ( n525 ) , ( n526 ) }  ;
assign n528 =  { ( n524 ) , ( n527 ) }  ;
assign n529 =  { ( n523 ) , ( n528 ) }  ;
assign n530 =  { ( n522 ) , ( n529 ) }  ;
assign n531 =  { ( n521 ) , ( n530 ) }  ;
assign n532 =  { ( n520 ) , ( n531 ) }  ;
assign n533 =  { ( n519 ) , ( n532 ) }  ;
assign n534 =  { ( n518 ) , ( n533 ) }  ;
assign n535 = n124[7:0] ;
assign n536 = LB2D_shift_7[7:0] ;
assign n537 = LB2D_shift_6[7:0] ;
assign n538 = LB2D_shift_5[7:0] ;
assign n539 = LB2D_shift_4[7:0] ;
assign n540 = LB2D_shift_3[7:0] ;
assign n541 = LB2D_shift_2[7:0] ;
assign n542 = LB2D_shift_1[7:0] ;
assign n543 = LB2D_shift_0[7:0] ;
assign n544 =  { ( n542 ) , ( n543 ) }  ;
assign n545 =  { ( n541 ) , ( n544 ) }  ;
assign n546 =  { ( n540 ) , ( n545 ) }  ;
assign n547 =  { ( n539 ) , ( n546 ) }  ;
assign n548 =  { ( n538 ) , ( n547 ) }  ;
assign n549 =  { ( n537 ) , ( n548 ) }  ;
assign n550 =  { ( n536 ) , ( n549 ) }  ;
assign n551 =  { ( n535 ) , ( n550 ) }  ;
assign n552 =  { ( n534 ) , ( n551 ) }  ;
assign n553 =  { ( n517 ) , ( n552 ) }  ;
assign n554 =  { ( n500 ) , ( n553 ) }  ;
assign n555 =  { ( n483 ) , ( n554 ) }  ;
assign n556 =  { ( n466 ) , ( n555 ) }  ;
assign n557 =  { ( n449 ) , ( n556 ) }  ;
assign n558 =  { ( n432 ) , ( n557 ) }  ;
assign n559 =  { ( n415 ) , ( n558 ) }  ;
assign n560 =  ( n398 ) ? ( n559 ) : ( stencil_stream_buff_0 ) ;
assign n561 =  ( n32 ) ? ( stencil_stream_buff_0 ) : ( stencil_stream_buff_0 ) ;
assign n562 =  ( n25 ) ? ( stencil_stream_buff_0 ) : ( n561 ) ;
assign n563 =  ( n20 ) ? ( n560 ) : ( n562 ) ;
assign n564 =  ( n13 ) ? ( stencil_stream_buff_0 ) : ( n563 ) ;
assign n565 =  ( n4 ) ? ( stencil_stream_buff_0 ) : ( n564 ) ;
assign n566 =  ( n32 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_1 ) ;
assign n567 =  ( n25 ) ? ( stencil_stream_buff_1 ) : ( n566 ) ;
assign n568 =  ( n20 ) ? ( stencil_stream_buff_0 ) : ( n567 ) ;
assign n569 =  ( n13 ) ? ( stencil_stream_buff_1 ) : ( n568 ) ;
assign n570 =  ( n4 ) ? ( stencil_stream_buff_1 ) : ( n569 ) ;
assign n571 =  ( n150 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n572 =  ( n18 ) ? ( stencil_stream_empty ) : ( 1'd0 ) ;
assign n573 =  ( n32 ) ? ( stencil_stream_empty ) : ( stencil_stream_empty ) ;
assign n574 =  ( n25 ) ? ( stencil_stream_empty ) : ( n573 ) ;
assign n575 =  ( n20 ) ? ( n572 ) : ( n574 ) ;
assign n576 =  ( n13 ) ? ( n571 ) : ( n575 ) ;
assign n577 =  ( n4 ) ? ( stencil_stream_empty ) : ( n576 ) ;
assign n578 =  ( n9 ) ? ( 1'd0 ) : ( 1'd0 ) ;
assign n579 =  ( stencil_stream_empty ) == ( 1'd1 )  ;
assign n580 =  ( n579 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n581 =  ( n18 ) ? ( stencil_stream_full ) : ( n580 ) ;
assign n582 =  ( n32 ) ? ( stencil_stream_full ) : ( stencil_stream_full ) ;
assign n583 =  ( n25 ) ? ( stencil_stream_full ) : ( n582 ) ;
assign n584 =  ( n20 ) ? ( n581 ) : ( n583 ) ;
assign n585 =  ( n13 ) ? ( n578 ) : ( n584 ) ;
assign n586 =  ( n4 ) ? ( stencil_stream_full ) : ( n585 ) ;
assign n587 = ~ ( n4 ) ;
assign n588 = ~ ( n13 ) ;
assign n589 =  ( n587 ) & ( n588 )  ;
assign n590 = ~ ( n20 ) ;
assign n591 =  ( n589 ) & ( n590 )  ;
assign n592 = ~ ( n25 ) ;
assign n593 =  ( n591 ) & ( n592 )  ;
assign n594 = ~ ( n32 ) ;
assign n595 =  ( n593 ) & ( n594 )  ;
assign n596 =  ( n593 ) & ( n32 )  ;
assign n597 =  ( n591 ) & ( n25 )  ;
assign n598 = ~ ( n291 ) ;
assign n599 =  ( n597 ) & ( n598 )  ;
assign n600 =  ( n597 ) & ( n291 )  ;
assign n601 =  ( n589 ) & ( n20 )  ;
assign n602 =  ( n587 ) & ( n13 )  ;
assign LB2D_proc_0_addr0 = n600 ? (n292) : (0);
assign LB2D_proc_0_data0 = n600 ? (n290) : (LB2D_proc_0[0]);
assign n603 = ~ ( n294 ) ;
assign n604 =  ( n597 ) & ( n603 )  ;
assign n605 =  ( n597 ) & ( n294 )  ;
assign LB2D_proc_1_addr0 = n605 ? (n292) : (0);
assign LB2D_proc_1_data0 = n605 ? (n290) : (LB2D_proc_1[0]);
assign n606 = ~ ( n296 ) ;
assign n607 =  ( n597 ) & ( n606 )  ;
assign n608 =  ( n597 ) & ( n296 )  ;
assign LB2D_proc_2_addr0 = n608 ? (n292) : (0);
assign LB2D_proc_2_data0 = n608 ? (n290) : (LB2D_proc_2[0]);
assign n609 = ~ ( n298 ) ;
assign n610 =  ( n597 ) & ( n609 )  ;
assign n611 =  ( n597 ) & ( n298 )  ;
assign LB2D_proc_3_addr0 = n611 ? (n292) : (0);
assign LB2D_proc_3_data0 = n611 ? (n290) : (LB2D_proc_3[0]);
assign n612 = ~ ( n300 ) ;
assign n613 =  ( n597 ) & ( n612 )  ;
assign n614 =  ( n597 ) & ( n300 )  ;
assign LB2D_proc_4_addr0 = n614 ? (n292) : (0);
assign LB2D_proc_4_data0 = n614 ? (n290) : (LB2D_proc_4[0]);
assign n615 = ~ ( n302 ) ;
assign n616 =  ( n597 ) & ( n615 )  ;
assign n617 =  ( n597 ) & ( n302 )  ;
assign LB2D_proc_5_addr0 = n617 ? (n292) : (0);
assign LB2D_proc_5_data0 = n617 ? (n290) : (LB2D_proc_5[0]);
assign n618 = ~ ( n304 ) ;
assign n619 =  ( n597 ) & ( n618 )  ;
assign n620 =  ( n597 ) & ( n304 )  ;
assign LB2D_proc_6_addr0 = n620 ? (n292) : (0);
assign LB2D_proc_6_data0 = n620 ? (n290) : (LB2D_proc_6[0]);
assign n621 = ~ ( n63 ) ;
assign n622 =  ( n597 ) & ( n621 )  ;
assign n623 =  ( n597 ) & ( n63 )  ;
assign LB2D_proc_7_addr0 = n623 ? (n292) : (0);
assign LB2D_proc_7_data0 = n623 ? (n290) : (LB2D_proc_7[0]);
/*
function [7:0] gb_fun ;
input [647:0] arg0;
    begin
//TODO: Add the specific function HERE.    end
endfunction
*/

always @(posedge clk) begin
   if(rst) begin
       LB1D_buff <= LB1D_buff;
       LB1D_in <= LB1D_in;
       LB1D_it_1 <= LB1D_it_1;
       LB1D_p_cnt <= LB1D_p_cnt;
       LB1D_uIn <= LB1D_uIn;
       LB2D_proc_w <= LB2D_proc_w;
       LB2D_proc_x <= LB2D_proc_x;
       LB2D_proc_y <= LB2D_proc_y;
       LB2D_shift_0 <= LB2D_shift_0;
       LB2D_shift_1 <= LB2D_shift_1;
       LB2D_shift_2 <= LB2D_shift_2;
       LB2D_shift_3 <= LB2D_shift_3;
       LB2D_shift_4 <= LB2D_shift_4;
       LB2D_shift_5 <= LB2D_shift_5;
       LB2D_shift_6 <= LB2D_shift_6;
       LB2D_shift_7 <= LB2D_shift_7;
       LB2D_shift_x <= LB2D_shift_x;
       LB2D_shift_y <= LB2D_shift_y;
       arg_0_TDATA <= arg_0_TDATA;
       arg_0_TVALID <= arg_0_TVALID;
       arg_1_TREADY <= arg_1_TREADY;
       gb_exit_it_1 <= gb_exit_it_1;
       gb_exit_it_2 <= gb_exit_it_2;
       gb_exit_it_3 <= gb_exit_it_3;
       gb_exit_it_4 <= gb_exit_it_4;
       gb_exit_it_5 <= gb_exit_it_5;
       gb_exit_it_6 <= gb_exit_it_6;
       gb_exit_it_7 <= gb_exit_it_7;
       gb_exit_it_8 <= gb_exit_it_8;
       gb_p_cnt <= gb_p_cnt;
       gb_pp_it_1 <= gb_pp_it_1;
       gb_pp_it_2 <= gb_pp_it_2;
       gb_pp_it_3 <= gb_pp_it_3;
       gb_pp_it_4 <= gb_pp_it_4;
       gb_pp_it_5 <= gb_pp_it_5;
       gb_pp_it_6 <= gb_pp_it_6;
       gb_pp_it_7 <= gb_pp_it_7;
       gb_pp_it_8 <= gb_pp_it_8;
       gb_pp_it_9 <= gb_pp_it_9;
       in_stream_buff_0 <= in_stream_buff_0;
       in_stream_buff_1 <= in_stream_buff_1;
       in_stream_empty <= in_stream_empty;
       in_stream_full <= in_stream_full;
       slice_stream_buff_0 <= slice_stream_buff_0;
       slice_stream_buff_1 <= slice_stream_buff_1;
       slice_stream_empty <= slice_stream_empty;
       slice_stream_full <= slice_stream_full;
       stencil_stream_buff_0 <= stencil_stream_buff_0;
       stencil_stream_buff_1 <= stencil_stream_buff_1;
       stencil_stream_empty <= stencil_stream_empty;
       stencil_stream_full <= stencil_stream_full;
   end
   else if(step) begin
       LB1D_buff <= n38;
       LB1D_in <= n44;
       LB1D_it_1 <= n45;
       LB1D_p_cnt <= n55;
       LB1D_uIn <= n61;
       LB2D_proc_w <= n71;
       LB2D_proc_x <= n78;
       LB2D_proc_y <= n87;
       LB2D_shift_0 <= n92;
       LB2D_shift_1 <= n97;
       LB2D_shift_2 <= n102;
       LB2D_shift_3 <= n107;
       LB2D_shift_4 <= n112;
       LB2D_shift_5 <= n117;
       LB2D_shift_6 <= n122;
       LB2D_shift_7 <= n129;
       LB2D_shift_x <= n139;
       LB2D_shift_y <= n149;
       arg_0_TDATA <= n157;
       arg_0_TVALID <= n164;
       arg_1_TREADY <= n170;
       gb_exit_it_1 <= n178;
       gb_exit_it_2 <= n183;
       gb_exit_it_3 <= n188;
       gb_exit_it_4 <= n193;
       gb_exit_it_5 <= n198;
       gb_exit_it_6 <= n203;
       gb_exit_it_7 <= n208;
       gb_exit_it_8 <= n213;
       gb_p_cnt <= n220;
       gb_pp_it_1 <= n225;
       gb_pp_it_2 <= n230;
       gb_pp_it_3 <= n235;
       gb_pp_it_4 <= n240;
       gb_pp_it_5 <= n245;
       gb_pp_it_6 <= n250;
       gb_pp_it_7 <= n255;
       gb_pp_it_8 <= n260;
       gb_pp_it_9 <= n265;
       in_stream_buff_0 <= n270;
       in_stream_buff_1 <= n275;
       in_stream_empty <= n282;
       in_stream_full <= n289;
       slice_stream_buff_0 <= n376;
       slice_stream_buff_1 <= n382;
       slice_stream_empty <= n389;
       slice_stream_full <= n397;
       stencil_stream_buff_0 <= n565;
       stencil_stream_buff_1 <= n570;
       stencil_stream_empty <= n577;
       stencil_stream_full <= n586;
       LB2D_proc_0 [ LB2D_proc_0_addr0 ] <= LB2D_proc_0_data0;
       LB2D_proc_1 [ LB2D_proc_1_addr0 ] <= LB2D_proc_1_data0;
       LB2D_proc_2 [ LB2D_proc_2_addr0 ] <= LB2D_proc_2_data0;
       LB2D_proc_3 [ LB2D_proc_3_addr0 ] <= LB2D_proc_3_data0;
       LB2D_proc_4 [ LB2D_proc_4_addr0 ] <= LB2D_proc_4_data0;
       LB2D_proc_5 [ LB2D_proc_5_addr0 ] <= LB2D_proc_5_data0;
       LB2D_proc_6 [ LB2D_proc_6_addr0 ] <= LB2D_proc_6_data0;
       LB2D_proc_7 [ LB2D_proc_7_addr0 ] <= LB2D_proc_7_data0;
   end
end
endmodule
