module GB(
arg_0_TREADY,
arg_1_TDATA,
arg_1_TVALID,
LB1D_buff,
LB1D_in,
LB1D_it_1,
LB1D_p_cnt,
LB2D_proc_w,
LB2D_proc_x,
LB2D_proc_y,
LB2D_shift_0,
LB2D_shift_1,
LB2D_shift_2,
LB2D_shift_3,
LB2D_shift_4,
LB2D_shift_5,
LB2D_shift_6,
LB2D_shift_7,
LB2D_shift_x,
LB2D_shift_y,
arg_0_TDATA,
arg_0_TVALID,
arg_1_TREADY,
gb_exit_it_1,
gb_exit_it_2,
gb_exit_it_3,
gb_exit_it_4,
gb_exit_it_5,
gb_exit_it_6,
gb_exit_it_7,
gb_exit_it_8,
gb_p_cnt,
gb_pp_it_1,
gb_pp_it_2,
gb_pp_it_3,
gb_pp_it_4,
gb_pp_it_5,
gb_pp_it_6,
gb_pp_it_7,
gb_pp_it_8,
gb_pp_it_9,
in_stream_buff_0,
in_stream_buff_1,
in_stream_empty,
in_stream_full,
slice_stream_buff_0,
slice_stream_buff_1,
slice_stream_empty,
slice_stream_full,
stencil_stream_buff_0,
stencil_stream_buff_1,
stencil_stream_empty,
stencil_stream_full,
clk,rst,
step
);
input            arg_0_TREADY;
input      [7:0] arg_1_TDATA;
input            arg_1_TVALID;
input clk;
input rst;
input step;
output      [7:0] LB1D_buff;
output      [7:0] LB1D_in;
output            LB1D_it_1;
output     [18:0] LB1D_p_cnt;
output     [63:0] LB2D_proc_w;
output      [8:0] LB2D_proc_x;
output      [9:0] LB2D_proc_y;
output     [71:0] LB2D_shift_0;
output     [71:0] LB2D_shift_1;
output     [71:0] LB2D_shift_2;
output     [71:0] LB2D_shift_3;
output     [71:0] LB2D_shift_4;
output     [71:0] LB2D_shift_5;
output     [71:0] LB2D_shift_6;
output     [71:0] LB2D_shift_7;
output      [8:0] LB2D_shift_x;
output      [9:0] LB2D_shift_y;
output      [7:0] arg_0_TDATA;
output            arg_0_TVALID;
output            arg_1_TREADY;
output            gb_exit_it_1;
output            gb_exit_it_2;
output            gb_exit_it_3;
output            gb_exit_it_4;
output            gb_exit_it_5;
output            gb_exit_it_6;
output            gb_exit_it_7;
output            gb_exit_it_8;
output     [18:0] gb_p_cnt;
output            gb_pp_it_1;
output            gb_pp_it_2;
output            gb_pp_it_3;
output            gb_pp_it_4;
output            gb_pp_it_5;
output            gb_pp_it_6;
output            gb_pp_it_7;
output            gb_pp_it_8;
output            gb_pp_it_9;
output      [7:0] in_stream_buff_0;
output      [7:0] in_stream_buff_1;
output            in_stream_empty;
output            in_stream_full;
output     [71:0] slice_stream_buff_0;
output     [71:0] slice_stream_buff_1;
output            slice_stream_empty;
output            slice_stream_full;
output    [647:0] stencil_stream_buff_0;
output    [647:0] stencil_stream_buff_1;
output            stencil_stream_empty;
output            stencil_stream_full;
reg      [7:0] LB1D_buff;
reg      [7:0] LB1D_in;
reg            LB1D_it_1;
reg     [18:0] LB1D_p_cnt;
reg     [63:0] LB2D_proc_w;
reg      [8:0] LB2D_proc_x;
reg      [9:0] LB2D_proc_y;
reg     [71:0] LB2D_shift_0;
reg     [71:0] LB2D_shift_1;
reg     [71:0] LB2D_shift_2;
reg     [71:0] LB2D_shift_3;
reg     [71:0] LB2D_shift_4;
reg     [71:0] LB2D_shift_5;
reg     [71:0] LB2D_shift_6;
reg     [71:0] LB2D_shift_7;
reg      [8:0] LB2D_shift_x;
reg      [9:0] LB2D_shift_y;
reg      [7:0] arg_0_TDATA;
reg            arg_0_TVALID;
reg            arg_1_TREADY;
reg            gb_exit_it_1;
reg            gb_exit_it_2;
reg            gb_exit_it_3;
reg            gb_exit_it_4;
reg            gb_exit_it_5;
reg            gb_exit_it_6;
reg            gb_exit_it_7;
reg            gb_exit_it_8;
reg     [18:0] gb_p_cnt;
reg            gb_pp_it_1;
reg            gb_pp_it_2;
reg            gb_pp_it_3;
reg            gb_pp_it_4;
reg            gb_pp_it_5;
reg            gb_pp_it_6;
reg            gb_pp_it_7;
reg            gb_pp_it_8;
reg            gb_pp_it_9;
reg      [7:0] in_stream_buff_0;
reg      [7:0] in_stream_buff_1;
reg            in_stream_empty;
reg            in_stream_full;
reg     [71:0] slice_stream_buff_0;
reg     [71:0] slice_stream_buff_1;
reg            slice_stream_empty;
reg            slice_stream_full;
reg    [647:0] stencil_stream_buff_0;
reg    [647:0] stencil_stream_buff_1;
reg            stencil_stream_empty;
reg            stencil_stream_full;
wire            arg_0_TREADY;
wire      [7:0] arg_1_TDATA;
wire            arg_1_TVALID;
wire            n0;
wire            n1;
wire            n2;
wire            n3;
wire            n4;
wire            n5;
wire            n6;
wire            n7;
wire            n8;
wire            n9;
wire            n10;
wire            n11;
wire            n12;
wire            n13;
wire            n14;
wire            n15;
wire            n16;
wire            n17;
wire            n18;
wire            n19;
wire            n20;
wire            n21;
wire            n22;
wire            n23;
wire            n24;
wire            n25;
wire            n26;
wire            n27;
wire            n28;
wire            n29;
wire            n30;
wire            n31;
wire            n32;
wire            n33;
wire            n34;
wire            n35;
wire            n36;
wire            n37;
wire      [7:0] n38;
wire      [7:0] n39;
wire      [7:0] n40;
wire      [7:0] n41;
wire      [7:0] n42;
wire      [7:0] n43;
wire      [7:0] n44;
wire      [7:0] n45;
wire      [7:0] n46;
wire      [7:0] n47;
wire      [7:0] n48;
wire            n49;
wire            n50;
wire            n51;
wire     [18:0] n52;
wire     [18:0] n53;
wire            n54;
wire     [18:0] n55;
wire     [18:0] n56;
wire     [18:0] n57;
wire     [18:0] n58;
wire     [18:0] n59;
wire     [18:0] n60;
wire     [18:0] n61;
wire     [18:0] n62;
wire            n63;
wire            n64;
wire     [63:0] n65;
wire     [63:0] n66;
wire     [63:0] n67;
wire     [63:0] n68;
wire     [63:0] n69;
wire     [63:0] n70;
wire     [63:0] n71;
wire     [63:0] n72;
wire     [63:0] n73;
wire            n74;
wire            n75;
wire            n76;
wire      [8:0] n77;
wire      [8:0] n78;
wire      [8:0] n79;
wire      [8:0] n80;
wire      [8:0] n81;
wire      [8:0] n82;
wire      [8:0] n83;
wire      [8:0] n84;
wire            n85;
wire      [9:0] n86;
wire      [9:0] n87;
wire      [9:0] n88;
wire      [9:0] n89;
wire      [9:0] n90;
wire      [9:0] n91;
wire      [9:0] n92;
wire            n93;
wire     [71:0] n94;
wire     [71:0] n95;
wire     [71:0] n96;
wire     [71:0] n97;
wire     [71:0] n98;
wire     [71:0] n99;
wire     [71:0] n100;
wire     [71:0] n101;
wire     [71:0] n102;
wire     [71:0] n103;
wire     [71:0] n104;
wire     [71:0] n105;
wire     [71:0] n106;
wire     [71:0] n107;
wire     [71:0] n108;
wire     [71:0] n109;
wire     [71:0] n110;
wire     [71:0] n111;
wire     [71:0] n112;
wire     [71:0] n113;
wire     [71:0] n114;
wire     [71:0] n115;
wire     [71:0] n116;
wire     [71:0] n117;
wire     [71:0] n118;
wire     [71:0] n119;
wire     [71:0] n120;
wire     [71:0] n121;
wire     [71:0] n122;
wire     [71:0] n123;
wire     [71:0] n124;
wire     [71:0] n125;
wire     [71:0] n126;
wire     [71:0] n127;
wire     [71:0] n128;
wire     [71:0] n129;
wire     [71:0] n130;
wire     [71:0] n131;
wire     [71:0] n132;
wire     [71:0] n133;
wire     [71:0] n134;
wire     [71:0] n135;
wire     [71:0] n136;
wire     [71:0] n137;
wire     [71:0] n138;
wire     [71:0] n139;
wire     [71:0] n140;
wire     [71:0] n141;
wire     [71:0] n142;
wire      [8:0] n143;
wire      [8:0] n144;
wire      [8:0] n145;
wire      [8:0] n146;
wire      [8:0] n147;
wire      [8:0] n148;
wire      [8:0] n149;
wire            n150;
wire            n151;
wire      [9:0] n152;
wire      [9:0] n153;
wire      [9:0] n154;
wire      [9:0] n155;
wire      [9:0] n156;
wire      [9:0] n157;
wire      [9:0] n158;
wire      [9:0] n159;
wire      [9:0] n160;
wire            n161;
wire    [647:0] n162;
wire      [7:0] n163;
wire      [7:0] n164;
wire      [7:0] n165;
wire      [7:0] n166;
wire      [7:0] n167;
wire      [7:0] n168;
wire      [7:0] n169;
wire            n170;
wire            n171;
wire            n172;
wire            n173;
wire            n174;
wire            n175;
wire            n176;
wire            n177;
wire            n178;
wire            n179;
wire            n180;
wire            n181;
wire            n182;
wire            n183;
wire            n184;
wire     [18:0] n185;
wire            n186;
wire            n187;
wire            n188;
wire            n189;
wire            n190;
wire            n191;
wire            n192;
wire            n193;
wire            n194;
wire            n195;
wire            n196;
wire            n197;
wire            n198;
wire            n199;
wire            n200;
wire            n201;
wire            n202;
wire            n203;
wire            n204;
wire            n205;
wire            n206;
wire            n207;
wire            n208;
wire            n209;
wire            n210;
wire            n211;
wire            n212;
wire            n213;
wire            n214;
wire            n215;
wire            n216;
wire            n217;
wire            n218;
wire            n219;
wire            n220;
wire            n221;
wire            n222;
wire            n223;
wire            n224;
wire            n225;
wire            n226;
wire            n227;
wire            n228;
wire            n229;
wire            n230;
wire            n231;
wire            n232;
wire            n233;
wire            n234;
wire            n235;
wire            n236;
wire     [18:0] n237;
wire     [18:0] n238;
wire     [18:0] n239;
wire     [18:0] n240;
wire     [18:0] n241;
wire     [18:0] n242;
wire     [18:0] n243;
wire            n244;
wire            n245;
wire            n246;
wire            n247;
wire            n248;
wire            n249;
wire            n250;
wire            n251;
wire            n252;
wire            n253;
wire            n254;
wire            n255;
wire            n256;
wire            n257;
wire            n258;
wire            n259;
wire            n260;
wire            n261;
wire            n262;
wire            n263;
wire            n264;
wire            n265;
wire            n266;
wire            n267;
wire            n268;
wire            n269;
wire            n270;
wire            n271;
wire            n272;
wire            n273;
wire            n274;
wire            n275;
wire            n276;
wire            n277;
wire            n278;
wire            n279;
wire            n280;
wire            n281;
wire            n282;
wire            n283;
wire            n284;
wire            n285;
wire            n286;
wire            n287;
wire            n288;
wire            n289;
wire            n290;
wire            n291;
wire            n292;
wire            n293;
wire            n294;
wire            n295;
wire            n296;
wire            n297;
wire      [7:0] n298;
wire      [7:0] n299;
wire      [7:0] n300;
wire      [7:0] n301;
wire      [7:0] n302;
wire      [7:0] n303;
wire      [7:0] n304;
wire      [7:0] n305;
wire      [7:0] n306;
wire      [7:0] n307;
wire      [7:0] n308;
wire      [7:0] n309;
wire            n310;
wire            n311;
wire            n312;
wire            n313;
wire            n314;
wire            n315;
wire            n316;
wire            n317;
wire            n318;
wire            n319;
wire            n320;
wire            n321;
wire            n322;
wire            n323;
wire            n324;
wire            n325;
wire      [7:0] n326;
wire            n327;
wire      [7:0] n328;
wire            n329;
wire      [7:0] n330;
wire            n331;
wire      [7:0] n332;
wire            n333;
wire      [7:0] n334;
wire            n335;
wire      [7:0] n336;
wire            n337;
wire      [7:0] n338;
wire            n339;
wire      [7:0] n340;
wire      [7:0] n341;
wire      [7:0] n342;
wire      [7:0] n343;
wire      [7:0] n344;
wire      [7:0] n345;
wire      [7:0] n346;
wire      [7:0] n347;
wire      [7:0] n348;
wire      [7:0] n349;
wire      [7:0] n350;
wire      [7:0] n351;
wire      [7:0] n352;
wire      [7:0] n353;
wire      [7:0] n354;
wire      [7:0] n355;
wire      [7:0] n356;
wire      [7:0] n357;
wire      [7:0] n358;
wire      [7:0] n359;
wire      [7:0] n360;
wire      [7:0] n361;
wire      [7:0] n362;
wire      [7:0] n363;
wire      [7:0] n364;
wire      [7:0] n365;
wire      [7:0] n366;
wire      [7:0] n367;
wire      [7:0] n368;
wire      [7:0] n369;
wire      [7:0] n370;
wire      [7:0] n371;
wire      [7:0] n372;
wire      [7:0] n373;
wire      [7:0] n374;
wire      [7:0] n375;
wire      [7:0] n376;
wire      [7:0] n377;
wire      [7:0] n378;
wire      [7:0] n379;
wire      [7:0] n380;
wire      [7:0] n381;
wire      [7:0] n382;
wire      [7:0] n383;
wire      [7:0] n384;
wire      [7:0] n385;
wire      [7:0] n386;
wire      [7:0] n387;
wire      [7:0] n388;
wire      [7:0] n389;
wire      [7:0] n390;
wire      [7:0] n391;
wire      [7:0] n392;
wire      [7:0] n393;
wire      [7:0] n394;
wire      [7:0] n395;
wire      [7:0] n396;
wire      [7:0] n397;
wire     [15:0] n398;
wire     [23:0] n399;
wire     [31:0] n400;
wire     [39:0] n401;
wire     [47:0] n402;
wire     [55:0] n403;
wire     [63:0] n404;
wire     [71:0] n405;
wire     [71:0] n406;
wire     [71:0] n407;
wire     [71:0] n408;
wire     [71:0] n409;
wire     [71:0] n410;
wire     [71:0] n411;
wire     [71:0] n412;
wire     [71:0] n413;
wire     [71:0] n414;
wire     [71:0] n415;
wire     [71:0] n416;
wire     [71:0] n417;
wire     [71:0] n418;
wire     [71:0] n419;
wire            n420;
wire            n421;
wire            n422;
wire            n423;
wire            n424;
wire            n425;
wire            n426;
wire            n427;
wire            n428;
wire            n429;
wire            n430;
wire            n431;
wire            n432;
wire            n433;
wire            n434;
wire            n435;
wire            n436;
wire            n437;
wire      [7:0] n438;
wire      [7:0] n439;
wire      [7:0] n440;
wire      [7:0] n441;
wire      [7:0] n442;
wire      [7:0] n443;
wire      [7:0] n444;
wire      [7:0] n445;
wire      [7:0] n446;
wire     [15:0] n447;
wire     [23:0] n448;
wire     [31:0] n449;
wire     [39:0] n450;
wire     [47:0] n451;
wire     [55:0] n452;
wire     [63:0] n453;
wire     [71:0] n454;
wire      [7:0] n455;
wire      [7:0] n456;
wire      [7:0] n457;
wire      [7:0] n458;
wire      [7:0] n459;
wire      [7:0] n460;
wire      [7:0] n461;
wire      [7:0] n462;
wire      [7:0] n463;
wire     [15:0] n464;
wire     [23:0] n465;
wire     [31:0] n466;
wire     [39:0] n467;
wire     [47:0] n468;
wire     [55:0] n469;
wire     [63:0] n470;
wire     [71:0] n471;
wire      [7:0] n472;
wire      [7:0] n473;
wire      [7:0] n474;
wire      [7:0] n475;
wire      [7:0] n476;
wire      [7:0] n477;
wire      [7:0] n478;
wire      [7:0] n479;
wire      [7:0] n480;
wire     [15:0] n481;
wire     [23:0] n482;
wire     [31:0] n483;
wire     [39:0] n484;
wire     [47:0] n485;
wire     [55:0] n486;
wire     [63:0] n487;
wire     [71:0] n488;
wire      [7:0] n489;
wire      [7:0] n490;
wire      [7:0] n491;
wire      [7:0] n492;
wire      [7:0] n493;
wire      [7:0] n494;
wire      [7:0] n495;
wire      [7:0] n496;
wire      [7:0] n497;
wire     [15:0] n498;
wire     [23:0] n499;
wire     [31:0] n500;
wire     [39:0] n501;
wire     [47:0] n502;
wire     [55:0] n503;
wire     [63:0] n504;
wire     [71:0] n505;
wire      [7:0] n506;
wire      [7:0] n507;
wire      [7:0] n508;
wire      [7:0] n509;
wire      [7:0] n510;
wire      [7:0] n511;
wire      [7:0] n512;
wire      [7:0] n513;
wire      [7:0] n514;
wire     [15:0] n515;
wire     [23:0] n516;
wire     [31:0] n517;
wire     [39:0] n518;
wire     [47:0] n519;
wire     [55:0] n520;
wire     [63:0] n521;
wire     [71:0] n522;
wire      [7:0] n523;
wire      [7:0] n524;
wire      [7:0] n525;
wire      [7:0] n526;
wire      [7:0] n527;
wire      [7:0] n528;
wire      [7:0] n529;
wire      [7:0] n530;
wire      [7:0] n531;
wire     [15:0] n532;
wire     [23:0] n533;
wire     [31:0] n534;
wire     [39:0] n535;
wire     [47:0] n536;
wire     [55:0] n537;
wire     [63:0] n538;
wire     [71:0] n539;
wire      [7:0] n540;
wire      [7:0] n541;
wire      [7:0] n542;
wire      [7:0] n543;
wire      [7:0] n544;
wire      [7:0] n545;
wire      [7:0] n546;
wire      [7:0] n547;
wire      [7:0] n548;
wire     [15:0] n549;
wire     [23:0] n550;
wire     [31:0] n551;
wire     [39:0] n552;
wire     [47:0] n553;
wire     [55:0] n554;
wire     [63:0] n555;
wire     [71:0] n556;
wire      [7:0] n557;
wire      [7:0] n558;
wire      [7:0] n559;
wire      [7:0] n560;
wire      [7:0] n561;
wire      [7:0] n562;
wire      [7:0] n563;
wire      [7:0] n564;
wire      [7:0] n565;
wire     [15:0] n566;
wire     [23:0] n567;
wire     [31:0] n568;
wire     [39:0] n569;
wire     [47:0] n570;
wire     [55:0] n571;
wire     [63:0] n572;
wire     [71:0] n573;
wire      [7:0] n574;
wire      [7:0] n575;
wire      [7:0] n576;
wire      [7:0] n577;
wire      [7:0] n578;
wire      [7:0] n579;
wire      [7:0] n580;
wire      [7:0] n581;
wire      [7:0] n582;
wire     [15:0] n583;
wire     [23:0] n584;
wire     [31:0] n585;
wire     [39:0] n586;
wire     [47:0] n587;
wire     [55:0] n588;
wire     [63:0] n589;
wire     [71:0] n590;
wire    [143:0] n591;
wire    [215:0] n592;
wire    [287:0] n593;
wire    [359:0] n594;
wire    [431:0] n595;
wire    [503:0] n596;
wire    [575:0] n597;
wire    [647:0] n598;
wire    [647:0] n599;
wire    [647:0] n600;
wire    [647:0] n601;
wire    [647:0] n602;
wire    [647:0] n603;
wire    [647:0] n604;
wire    [647:0] n605;
wire    [647:0] n606;
wire    [647:0] n607;
wire    [647:0] n608;
wire    [647:0] n609;
wire    [647:0] n610;
wire    [647:0] n611;
wire            n612;
wire            n613;
wire            n614;
wire            n615;
wire            n616;
wire            n617;
wire            n618;
wire            n619;
wire            n620;
wire            n621;
wire            n622;
wire            n623;
wire            n624;
wire            n625;
wire            n626;
wire            n627;
wire            n628;
wire            n629;
wire      [8:0] LB2D_proc_0_addr0;
wire      [7:0] LB2D_proc_0_data0;
wire            n630;
wire            n631;
wire            n632;
wire            n633;
wire            n634;
wire            n635;
wire            n636;
wire            n637;
wire            n638;
wire            n639;
wire            n640;
wire            n641;
wire            n642;
wire            n643;
wire            n644;
wire            n645;
wire            n646;
wire            n647;
wire            n648;
wire      [8:0] LB2D_proc_1_addr0;
wire      [7:0] LB2D_proc_1_data0;
wire            n649;
wire            n650;
wire            n651;
wire      [8:0] LB2D_proc_2_addr0;
wire      [7:0] LB2D_proc_2_data0;
wire            n652;
wire            n653;
wire            n654;
wire      [8:0] LB2D_proc_3_addr0;
wire      [7:0] LB2D_proc_3_data0;
wire            n655;
wire            n656;
wire            n657;
wire      [8:0] LB2D_proc_4_addr0;
wire      [7:0] LB2D_proc_4_data0;
wire            n658;
wire            n659;
wire            n660;
wire      [8:0] LB2D_proc_5_addr0;
wire      [7:0] LB2D_proc_5_data0;
wire            n661;
wire            n662;
wire            n663;
wire      [8:0] LB2D_proc_6_addr0;
wire      [7:0] LB2D_proc_6_data0;
wire            n664;
wire            n665;
wire            n666;
wire      [8:0] LB2D_proc_7_addr0;
wire      [7:0] LB2D_proc_7_data0;
wire            n667;
wire            n668;
wire            n669;
wire            n670;
reg      [7:0] LB2D_proc_0[511:0];
reg      [7:0] LB2D_proc_1[511:0];
reg      [7:0] LB2D_proc_2[511:0];
reg      [7:0] LB2D_proc_3[511:0];
reg      [7:0] LB2D_proc_4[511:0];
reg      [7:0] LB2D_proc_5[511:0];
reg      [7:0] LB2D_proc_6[511:0];
reg      [7:0] LB2D_proc_7[511:0];
wire clk;
wire rst;
wire step;
assign n0 =  ( arg_0_TREADY ) == ( 1'd1 )  ;
assign n1 =  ( arg_0_TVALID ) == ( 1'd1 )  ;
assign n2 =  ( n0 ) & ( n1 )  ;
assign n3 =  ( arg_1_TVALID ) == ( 1'd0 )  ;
assign n4 =  ( n2 ) & ( n3 )  ;
assign n5 =  ( arg_1_TREADY ) == ( 1'd1 )  ;
assign n6 =  ( arg_1_TVALID ) == ( 1'd1 )  ;
assign n7 =  ( n5 ) & ( n6 )  ;
assign n8 =  ( arg_0_TREADY ) == ( 1'd0 )  ;
assign n9 =  ( n7 ) & ( n8 )  ;
assign n10 =  ( arg_0_TVALID ) == ( 1'd0 )  ;
assign n11 =  ( gb_exit_it_1 ) == ( 1'd0 )  ;
assign n12 =  ( stencil_stream_empty ) == ( 1'd0 )  ;
assign n13 =  ( n11 ) & ( n12 )  ;
assign n14 =  ( gb_exit_it_1 ) == ( 1'd1 )  ;
assign n15 =  ( gb_exit_it_8 ) == ( 1'd0 )  ;
assign n16 =  ( n14 ) & ( n15 )  ;
assign n17 =  ( n13 ) | ( n16 )  ;
assign n18 =  ( n10 ) & ( n17 )  ;
assign n19 =  ( slice_stream_empty ) == ( 1'd0 )  ;
assign n20 =  ( LB2D_shift_x ) != ( 9'd488 )  ;
assign n21 =  ( n19 ) & ( n20 )  ;
assign n22 =  ( stencil_stream_full ) == ( 1'd0 )  ;
assign n23 =  ( LB2D_shift_x ) < ( 9'd8 )  ;
assign n24 =  ( n22 ) | ( n23 )  ;
assign n25 =  ( n21 ) & ( n24 )  ;
assign n26 =  ( in_stream_empty ) == ( 1'd0 )  ;
assign n27 =  ( LB2D_proc_x ) != ( 9'd488 )  ;
assign n28 =  ( n26 ) & ( n27 )  ;
assign n29 =  ( slice_stream_full ) == ( 1'd0 )  ;
assign n30 =  ( LB2D_proc_y ) < ( 10'd8 )  ;
assign n31 =  ( n29 ) | ( n30 )  ;
assign n32 =  ( n28 ) & ( n31 )  ;
assign n33 =  ( arg_1_TREADY ) == ( 1'd0 )  ;
assign n34 =  ( in_stream_full ) == ( 1'd0 )  ;
assign n35 =  ( n33 ) & ( n34 )  ;
assign n36 =  ( LB1D_it_1 ) == ( 1'd1 )  ;
assign n37 =  ( n35 ) & ( n36 )  ;
assign n38 =  ( n37 ) ? ( LB1D_in ) : ( LB1D_buff ) ;
assign n39 =  ( n32 ) ? ( LB1D_buff ) : ( n38 ) ;
assign n40 =  ( n25 ) ? ( LB1D_buff ) : ( n39 ) ;
assign n41 =  ( n18 ) ? ( LB1D_buff ) : ( n40 ) ;
assign n42 =  ( n9 ) ? ( LB1D_buff ) : ( n41 ) ;
assign n43 =  ( n4 ) ? ( LB1D_buff ) : ( n42 ) ;
assign n44 =  ( n37 ) ? ( arg_1_TDATA ) : ( LB1D_in ) ;
assign n45 =  ( n25 ) ? ( LB1D_in ) : ( n44 ) ;
assign n46 =  ( n18 ) ? ( LB1D_in ) : ( n45 ) ;
assign n47 =  ( n9 ) ? ( LB1D_in ) : ( n46 ) ;
assign n48 =  ( n4 ) ? ( LB1D_in ) : ( n47 ) ;
assign n49 =  ( LB1D_it_1 ) == ( 1'd0 )  ;
assign n50 =  ( n35 ) & ( n49 )  ;
assign n51 =  ( n50 ) ? ( 1'd1 ) : ( LB1D_it_1 ) ;
assign n52 =  ( LB1D_p_cnt ) + ( 19'd1 )  ;
assign n53 =  ( 19'd316224 ) - ( 19'd1 )  ;
assign n54 =  ( LB1D_p_cnt ) == ( n53 )  ;
assign n55 =  ( n54 ) ? ( 19'd0 ) : ( n52 ) ;
assign n56 =  ( n37 ) ? ( n55 ) : ( LB1D_p_cnt ) ;
assign n57 =  ( n50 ) ? ( n52 ) : ( n56 ) ;
assign n58 =  ( n32 ) ? ( LB1D_p_cnt ) : ( n57 ) ;
assign n59 =  ( n25 ) ? ( LB1D_p_cnt ) : ( n58 ) ;
assign n60 =  ( n18 ) ? ( LB1D_p_cnt ) : ( n59 ) ;
assign n61 =  ( n9 ) ? ( LB1D_p_cnt ) : ( n60 ) ;
assign n62 =  ( n4 ) ? ( LB1D_p_cnt ) : ( n61 ) ;
assign n63 =  ( LB2D_proc_w ) < ( 64'd7 )  ;
assign n64 =  ( LB2D_proc_x ) < ( 9'd488 )  ;
assign n65 =  ( LB2D_proc_w ) + ( 64'd1 )  ;
assign n66 =  ( n64 ) ? ( LB2D_proc_w ) : ( n65 ) ;
assign n67 =  ( n63 ) ? ( n66 ) : ( 64'd0 ) ;
assign n68 =  ( n37 ) ? ( LB2D_proc_w ) : ( LB2D_proc_w ) ;
assign n69 =  ( n32 ) ? ( n67 ) : ( n68 ) ;
assign n70 =  ( n25 ) ? ( LB2D_proc_w ) : ( n69 ) ;
assign n71 =  ( n18 ) ? ( LB2D_proc_w ) : ( n70 ) ;
assign n72 =  ( n9 ) ? ( LB2D_proc_w ) : ( n71 ) ;
assign n73 =  ( n4 ) ? ( LB2D_proc_w ) : ( n72 ) ;
assign n74 =  ( LB2D_proc_x ) == ( 9'd488 )  ;
assign n75 =  ( n26 ) & ( n74 )  ;
assign n76 =  ( n75 ) & ( n31 )  ;
assign n77 =  ( LB2D_proc_x ) + ( 9'd1 )  ;
assign n78 =  ( n37 ) ? ( LB2D_proc_x ) : ( LB2D_proc_x ) ;
assign n79 =  ( n32 ) ? ( n77 ) : ( n78 ) ;
assign n80 =  ( n76 ) ? ( 9'd0 ) : ( n79 ) ;
assign n81 =  ( n25 ) ? ( LB2D_proc_x ) : ( n80 ) ;
assign n82 =  ( n18 ) ? ( LB2D_proc_x ) : ( n81 ) ;
assign n83 =  ( n9 ) ? ( LB2D_proc_x ) : ( n82 ) ;
assign n84 =  ( n4 ) ? ( LB2D_proc_x ) : ( n83 ) ;
assign n85 =  ( LB2D_proc_y ) < ( 10'd488 )  ;
assign n86 =  ( n85 ) ? ( LB2D_proc_y ) : ( 10'd488 ) ;
assign n87 =  ( n37 ) ? ( LB2D_proc_y ) : ( LB2D_proc_y ) ;
assign n88 =  ( n32 ) ? ( n86 ) : ( n87 ) ;
assign n89 =  ( n25 ) ? ( LB2D_proc_y ) : ( n88 ) ;
assign n90 =  ( n18 ) ? ( LB2D_proc_y ) : ( n89 ) ;
assign n91 =  ( n9 ) ? ( LB2D_proc_y ) : ( n90 ) ;
assign n92 =  ( n4 ) ? ( LB2D_proc_y ) : ( n91 ) ;
assign n93 =  ( slice_stream_full ) == ( 1'd1 )  ;
assign n94 =  ( n93 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n95 =  ( n37 ) ? ( LB2D_shift_0 ) : ( LB2D_shift_0 ) ;
assign n96 =  ( n32 ) ? ( LB2D_shift_0 ) : ( n95 ) ;
assign n97 =  ( n25 ) ? ( n94 ) : ( n96 ) ;
assign n98 =  ( n18 ) ? ( LB2D_shift_0 ) : ( n97 ) ;
assign n99 =  ( n9 ) ? ( LB2D_shift_0 ) : ( n98 ) ;
assign n100 =  ( n4 ) ? ( LB2D_shift_0 ) : ( n99 ) ;
assign n101 =  ( n37 ) ? ( LB2D_shift_1 ) : ( LB2D_shift_1 ) ;
assign n102 =  ( n32 ) ? ( LB2D_shift_1 ) : ( n101 ) ;
assign n103 =  ( n25 ) ? ( LB2D_shift_0 ) : ( n102 ) ;
assign n104 =  ( n18 ) ? ( LB2D_shift_1 ) : ( n103 ) ;
assign n105 =  ( n9 ) ? ( LB2D_shift_1 ) : ( n104 ) ;
assign n106 =  ( n4 ) ? ( LB2D_shift_1 ) : ( n105 ) ;
assign n107 =  ( n37 ) ? ( LB2D_shift_2 ) : ( LB2D_shift_2 ) ;
assign n108 =  ( n32 ) ? ( LB2D_shift_2 ) : ( n107 ) ;
assign n109 =  ( n25 ) ? ( LB2D_shift_1 ) : ( n108 ) ;
assign n110 =  ( n18 ) ? ( LB2D_shift_2 ) : ( n109 ) ;
assign n111 =  ( n9 ) ? ( LB2D_shift_2 ) : ( n110 ) ;
assign n112 =  ( n4 ) ? ( LB2D_shift_2 ) : ( n111 ) ;
assign n113 =  ( n37 ) ? ( LB2D_shift_3 ) : ( LB2D_shift_3 ) ;
assign n114 =  ( n32 ) ? ( LB2D_shift_3 ) : ( n113 ) ;
assign n115 =  ( n25 ) ? ( LB2D_shift_2 ) : ( n114 ) ;
assign n116 =  ( n18 ) ? ( LB2D_shift_3 ) : ( n115 ) ;
assign n117 =  ( n9 ) ? ( LB2D_shift_3 ) : ( n116 ) ;
assign n118 =  ( n4 ) ? ( LB2D_shift_3 ) : ( n117 ) ;
assign n119 =  ( n37 ) ? ( LB2D_shift_4 ) : ( LB2D_shift_4 ) ;
assign n120 =  ( n32 ) ? ( LB2D_shift_4 ) : ( n119 ) ;
assign n121 =  ( n25 ) ? ( LB2D_shift_3 ) : ( n120 ) ;
assign n122 =  ( n18 ) ? ( LB2D_shift_4 ) : ( n121 ) ;
assign n123 =  ( n9 ) ? ( LB2D_shift_4 ) : ( n122 ) ;
assign n124 =  ( n4 ) ? ( LB2D_shift_4 ) : ( n123 ) ;
assign n125 =  ( n37 ) ? ( LB2D_shift_5 ) : ( LB2D_shift_5 ) ;
assign n126 =  ( n32 ) ? ( LB2D_shift_5 ) : ( n125 ) ;
assign n127 =  ( n25 ) ? ( LB2D_shift_4 ) : ( n126 ) ;
assign n128 =  ( n18 ) ? ( LB2D_shift_5 ) : ( n127 ) ;
assign n129 =  ( n9 ) ? ( LB2D_shift_5 ) : ( n128 ) ;
assign n130 =  ( n4 ) ? ( LB2D_shift_5 ) : ( n129 ) ;
assign n131 =  ( n37 ) ? ( LB2D_shift_6 ) : ( LB2D_shift_6 ) ;
assign n132 =  ( n32 ) ? ( LB2D_shift_6 ) : ( n131 ) ;
assign n133 =  ( n25 ) ? ( LB2D_shift_5 ) : ( n132 ) ;
assign n134 =  ( n18 ) ? ( LB2D_shift_6 ) : ( n133 ) ;
assign n135 =  ( n9 ) ? ( LB2D_shift_6 ) : ( n134 ) ;
assign n136 =  ( n4 ) ? ( LB2D_shift_6 ) : ( n135 ) ;
assign n137 =  ( n37 ) ? ( LB2D_shift_7 ) : ( LB2D_shift_7 ) ;
assign n138 =  ( n32 ) ? ( LB2D_shift_7 ) : ( n137 ) ;
assign n139 =  ( n25 ) ? ( LB2D_shift_6 ) : ( n138 ) ;
assign n140 =  ( n18 ) ? ( LB2D_shift_7 ) : ( n139 ) ;
assign n141 =  ( n9 ) ? ( LB2D_shift_7 ) : ( n140 ) ;
assign n142 =  ( n4 ) ? ( LB2D_shift_7 ) : ( n141 ) ;
assign n143 =  ( LB2D_shift_x ) + ( 9'd1 )  ;
assign n144 =  ( n37 ) ? ( LB2D_shift_x ) : ( LB2D_shift_x ) ;
assign n145 =  ( n32 ) ? ( LB2D_shift_x ) : ( n144 ) ;
assign n146 =  ( n25 ) ? ( n143 ) : ( n145 ) ;
assign n147 =  ( n18 ) ? ( LB2D_shift_x ) : ( n146 ) ;
assign n148 =  ( n9 ) ? ( LB2D_shift_x ) : ( n147 ) ;
assign n149 =  ( n4 ) ? ( LB2D_shift_x ) : ( n148 ) ;
assign n150 =  ( LB2D_shift_y ) < ( 10'd480 )  ;
assign n151 =  ( LB2D_shift_x ) < ( 9'd488 )  ;
assign n152 =  ( LB2D_shift_y ) + ( 10'd1 )  ;
assign n153 =  ( n151 ) ? ( LB2D_shift_y ) : ( n152 ) ;
assign n154 =  ( n150 ) ? ( n153 ) : ( 10'd480 ) ;
assign n155 =  ( n37 ) ? ( LB2D_shift_y ) : ( LB2D_shift_y ) ;
assign n156 =  ( n32 ) ? ( LB2D_shift_y ) : ( n155 ) ;
assign n157 =  ( n25 ) ? ( n154 ) : ( n156 ) ;
assign n158 =  ( n18 ) ? ( LB2D_shift_y ) : ( n157 ) ;
assign n159 =  ( n9 ) ? ( LB2D_shift_y ) : ( n158 ) ;
assign n160 =  ( n4 ) ? ( LB2D_shift_y ) : ( n159 ) ;
assign n161 =  ( stencil_stream_full ) == ( 1'd1 )  ;
assign n162 =  ( n161 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_0 ) ;
assign n163 = gb_fun(n162) ;
assign n164 =  ( n37 ) ? ( arg_0_TDATA ) : ( arg_0_TDATA ) ;
assign n165 =  ( n32 ) ? ( arg_0_TDATA ) : ( n164 ) ;
assign n166 =  ( n25 ) ? ( arg_0_TDATA ) : ( n165 ) ;
assign n167 =  ( n18 ) ? ( n163 ) : ( n166 ) ;
assign n168 =  ( n9 ) ? ( arg_0_TDATA ) : ( n167 ) ;
assign n169 =  ( n4 ) ? ( arg_0_TDATA ) : ( n168 ) ;
assign n170 =  ( gb_pp_it_8 ) == ( 1'd1 )  ;
assign n171 =  ( n170 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n172 =  ( n37 ) ? ( arg_0_TVALID ) : ( arg_0_TVALID ) ;
assign n173 =  ( n32 ) ? ( arg_0_TVALID ) : ( n172 ) ;
assign n174 =  ( n25 ) ? ( arg_0_TVALID ) : ( n173 ) ;
assign n175 =  ( n18 ) ? ( n171 ) : ( n174 ) ;
assign n176 =  ( n9 ) ? ( arg_0_TVALID ) : ( n175 ) ;
assign n177 =  ( n4 ) ? ( 1'd0 ) : ( n176 ) ;
assign n178 =  ( n37 ) ? ( 1'd1 ) : ( arg_1_TREADY ) ;
assign n179 =  ( n50 ) ? ( 1'd1 ) : ( n178 ) ;
assign n180 =  ( n32 ) ? ( arg_1_TREADY ) : ( n179 ) ;
assign n181 =  ( n25 ) ? ( arg_1_TREADY ) : ( n180 ) ;
assign n182 =  ( n18 ) ? ( arg_1_TREADY ) : ( n181 ) ;
assign n183 =  ( n9 ) ? ( 1'd0 ) : ( n182 ) ;
assign n184 =  ( n4 ) ? ( 1'd0 ) : ( n183 ) ;
assign n185 =  ( gb_p_cnt ) + ( 19'd1 )  ;
assign n186 =  ( n185 ) == ( 19'd307200 )  ;
assign n187 =  ( n186 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n188 =  ( n37 ) ? ( gb_exit_it_1 ) : ( gb_exit_it_1 ) ;
assign n189 =  ( n32 ) ? ( gb_exit_it_1 ) : ( n188 ) ;
assign n190 =  ( n25 ) ? ( gb_exit_it_1 ) : ( n189 ) ;
assign n191 =  ( n18 ) ? ( n187 ) : ( n190 ) ;
assign n192 =  ( n9 ) ? ( gb_exit_it_1 ) : ( n191 ) ;
assign n193 =  ( n4 ) ? ( gb_exit_it_1 ) : ( n192 ) ;
assign n194 =  ( n37 ) ? ( gb_exit_it_2 ) : ( gb_exit_it_2 ) ;
assign n195 =  ( n32 ) ? ( gb_exit_it_2 ) : ( n194 ) ;
assign n196 =  ( n25 ) ? ( gb_exit_it_2 ) : ( n195 ) ;
assign n197 =  ( n18 ) ? ( gb_exit_it_1 ) : ( n196 ) ;
assign n198 =  ( n9 ) ? ( gb_exit_it_2 ) : ( n197 ) ;
assign n199 =  ( n4 ) ? ( gb_exit_it_2 ) : ( n198 ) ;
assign n200 =  ( n37 ) ? ( gb_exit_it_3 ) : ( gb_exit_it_3 ) ;
assign n201 =  ( n32 ) ? ( gb_exit_it_3 ) : ( n200 ) ;
assign n202 =  ( n25 ) ? ( gb_exit_it_3 ) : ( n201 ) ;
assign n203 =  ( n18 ) ? ( gb_exit_it_2 ) : ( n202 ) ;
assign n204 =  ( n9 ) ? ( gb_exit_it_3 ) : ( n203 ) ;
assign n205 =  ( n4 ) ? ( gb_exit_it_3 ) : ( n204 ) ;
assign n206 =  ( n37 ) ? ( gb_exit_it_4 ) : ( gb_exit_it_4 ) ;
assign n207 =  ( n32 ) ? ( gb_exit_it_4 ) : ( n206 ) ;
assign n208 =  ( n25 ) ? ( gb_exit_it_4 ) : ( n207 ) ;
assign n209 =  ( n18 ) ? ( gb_exit_it_3 ) : ( n208 ) ;
assign n210 =  ( n9 ) ? ( gb_exit_it_4 ) : ( n209 ) ;
assign n211 =  ( n4 ) ? ( gb_exit_it_4 ) : ( n210 ) ;
assign n212 =  ( n37 ) ? ( gb_exit_it_5 ) : ( gb_exit_it_5 ) ;
assign n213 =  ( n32 ) ? ( gb_exit_it_5 ) : ( n212 ) ;
assign n214 =  ( n25 ) ? ( gb_exit_it_5 ) : ( n213 ) ;
assign n215 =  ( n18 ) ? ( gb_exit_it_4 ) : ( n214 ) ;
assign n216 =  ( n9 ) ? ( gb_exit_it_5 ) : ( n215 ) ;
assign n217 =  ( n4 ) ? ( gb_exit_it_5 ) : ( n216 ) ;
assign n218 =  ( n37 ) ? ( gb_exit_it_6 ) : ( gb_exit_it_6 ) ;
assign n219 =  ( n32 ) ? ( gb_exit_it_6 ) : ( n218 ) ;
assign n220 =  ( n25 ) ? ( gb_exit_it_6 ) : ( n219 ) ;
assign n221 =  ( n18 ) ? ( gb_exit_it_5 ) : ( n220 ) ;
assign n222 =  ( n9 ) ? ( gb_exit_it_6 ) : ( n221 ) ;
assign n223 =  ( n4 ) ? ( gb_exit_it_6 ) : ( n222 ) ;
assign n224 =  ( n37 ) ? ( gb_exit_it_7 ) : ( gb_exit_it_7 ) ;
assign n225 =  ( n32 ) ? ( gb_exit_it_7 ) : ( n224 ) ;
assign n226 =  ( n25 ) ? ( gb_exit_it_7 ) : ( n225 ) ;
assign n227 =  ( n18 ) ? ( gb_exit_it_6 ) : ( n226 ) ;
assign n228 =  ( n9 ) ? ( gb_exit_it_7 ) : ( n227 ) ;
assign n229 =  ( n4 ) ? ( gb_exit_it_7 ) : ( n228 ) ;
assign n230 =  ( n37 ) ? ( gb_exit_it_8 ) : ( gb_exit_it_8 ) ;
assign n231 =  ( n32 ) ? ( gb_exit_it_8 ) : ( n230 ) ;
assign n232 =  ( n25 ) ? ( gb_exit_it_8 ) : ( n231 ) ;
assign n233 =  ( n18 ) ? ( gb_exit_it_7 ) : ( n232 ) ;
assign n234 =  ( n9 ) ? ( gb_exit_it_8 ) : ( n233 ) ;
assign n235 =  ( n4 ) ? ( gb_exit_it_8 ) : ( n234 ) ;
assign n236 =  ( gb_p_cnt ) < ( 19'd307200 )  ;
assign n237 =  ( n236 ) ? ( n185 ) : ( 19'd307200 ) ;
assign n238 =  ( n37 ) ? ( gb_p_cnt ) : ( gb_p_cnt ) ;
assign n239 =  ( n32 ) ? ( gb_p_cnt ) : ( n238 ) ;
assign n240 =  ( n25 ) ? ( gb_p_cnt ) : ( n239 ) ;
assign n241 =  ( n18 ) ? ( n237 ) : ( n240 ) ;
assign n242 =  ( n9 ) ? ( gb_p_cnt ) : ( n241 ) ;
assign n243 =  ( n4 ) ? ( gb_p_cnt ) : ( n242 ) ;
assign n244 =  ( n37 ) ? ( gb_pp_it_1 ) : ( gb_pp_it_1 ) ;
assign n245 =  ( n32 ) ? ( gb_pp_it_1 ) : ( n244 ) ;
assign n246 =  ( n25 ) ? ( gb_pp_it_1 ) : ( n245 ) ;
assign n247 =  ( n18 ) ? ( 1'd1 ) : ( n246 ) ;
assign n248 =  ( n9 ) ? ( gb_pp_it_1 ) : ( n247 ) ;
assign n249 =  ( n4 ) ? ( gb_pp_it_1 ) : ( n248 ) ;
assign n250 =  ( n37 ) ? ( gb_pp_it_2 ) : ( gb_pp_it_2 ) ;
assign n251 =  ( n32 ) ? ( gb_pp_it_2 ) : ( n250 ) ;
assign n252 =  ( n25 ) ? ( gb_pp_it_2 ) : ( n251 ) ;
assign n253 =  ( n18 ) ? ( gb_pp_it_1 ) : ( n252 ) ;
assign n254 =  ( n9 ) ? ( gb_pp_it_2 ) : ( n253 ) ;
assign n255 =  ( n4 ) ? ( gb_pp_it_2 ) : ( n254 ) ;
assign n256 =  ( n37 ) ? ( gb_pp_it_3 ) : ( gb_pp_it_3 ) ;
assign n257 =  ( n32 ) ? ( gb_pp_it_3 ) : ( n256 ) ;
assign n258 =  ( n25 ) ? ( gb_pp_it_3 ) : ( n257 ) ;
assign n259 =  ( n18 ) ? ( gb_pp_it_2 ) : ( n258 ) ;
assign n260 =  ( n9 ) ? ( gb_pp_it_3 ) : ( n259 ) ;
assign n261 =  ( n4 ) ? ( gb_pp_it_3 ) : ( n260 ) ;
assign n262 =  ( n37 ) ? ( gb_pp_it_4 ) : ( gb_pp_it_4 ) ;
assign n263 =  ( n32 ) ? ( gb_pp_it_4 ) : ( n262 ) ;
assign n264 =  ( n25 ) ? ( gb_pp_it_4 ) : ( n263 ) ;
assign n265 =  ( n18 ) ? ( gb_pp_it_3 ) : ( n264 ) ;
assign n266 =  ( n9 ) ? ( gb_pp_it_4 ) : ( n265 ) ;
assign n267 =  ( n4 ) ? ( gb_pp_it_4 ) : ( n266 ) ;
assign n268 =  ( n37 ) ? ( gb_pp_it_5 ) : ( gb_pp_it_5 ) ;
assign n269 =  ( n32 ) ? ( gb_pp_it_5 ) : ( n268 ) ;
assign n270 =  ( n25 ) ? ( gb_pp_it_5 ) : ( n269 ) ;
assign n271 =  ( n18 ) ? ( gb_pp_it_4 ) : ( n270 ) ;
assign n272 =  ( n9 ) ? ( gb_pp_it_5 ) : ( n271 ) ;
assign n273 =  ( n4 ) ? ( gb_pp_it_5 ) : ( n272 ) ;
assign n274 =  ( n37 ) ? ( gb_pp_it_6 ) : ( gb_pp_it_6 ) ;
assign n275 =  ( n32 ) ? ( gb_pp_it_6 ) : ( n274 ) ;
assign n276 =  ( n25 ) ? ( gb_pp_it_6 ) : ( n275 ) ;
assign n277 =  ( n18 ) ? ( gb_pp_it_5 ) : ( n276 ) ;
assign n278 =  ( n9 ) ? ( gb_pp_it_6 ) : ( n277 ) ;
assign n279 =  ( n4 ) ? ( gb_pp_it_6 ) : ( n278 ) ;
assign n280 =  ( n37 ) ? ( gb_pp_it_7 ) : ( gb_pp_it_7 ) ;
assign n281 =  ( n32 ) ? ( gb_pp_it_7 ) : ( n280 ) ;
assign n282 =  ( n25 ) ? ( gb_pp_it_7 ) : ( n281 ) ;
assign n283 =  ( n18 ) ? ( gb_pp_it_6 ) : ( n282 ) ;
assign n284 =  ( n9 ) ? ( gb_pp_it_7 ) : ( n283 ) ;
assign n285 =  ( n4 ) ? ( gb_pp_it_7 ) : ( n284 ) ;
assign n286 =  ( n37 ) ? ( gb_pp_it_8 ) : ( gb_pp_it_8 ) ;
assign n287 =  ( n32 ) ? ( gb_pp_it_8 ) : ( n286 ) ;
assign n288 =  ( n25 ) ? ( gb_pp_it_8 ) : ( n287 ) ;
assign n289 =  ( n18 ) ? ( gb_pp_it_7 ) : ( n288 ) ;
assign n290 =  ( n9 ) ? ( gb_pp_it_8 ) : ( n289 ) ;
assign n291 =  ( n4 ) ? ( gb_pp_it_8 ) : ( n290 ) ;
assign n292 =  ( n37 ) ? ( gb_pp_it_9 ) : ( gb_pp_it_9 ) ;
assign n293 =  ( n32 ) ? ( gb_pp_it_9 ) : ( n292 ) ;
assign n294 =  ( n25 ) ? ( gb_pp_it_9 ) : ( n293 ) ;
assign n295 =  ( n18 ) ? ( gb_pp_it_8 ) : ( n294 ) ;
assign n296 =  ( n9 ) ? ( gb_pp_it_9 ) : ( n295 ) ;
assign n297 =  ( n4 ) ? ( gb_pp_it_9 ) : ( n296 ) ;
assign n298 =  ( n37 ) ? ( LB1D_buff ) : ( in_stream_buff_0 ) ;
assign n299 =  ( n32 ) ? ( in_stream_buff_0 ) : ( n298 ) ;
assign n300 =  ( n25 ) ? ( in_stream_buff_0 ) : ( n299 ) ;
assign n301 =  ( n18 ) ? ( in_stream_buff_0 ) : ( n300 ) ;
assign n302 =  ( n9 ) ? ( in_stream_buff_0 ) : ( n301 ) ;
assign n303 =  ( n4 ) ? ( in_stream_buff_0 ) : ( n302 ) ;
assign n304 =  ( n37 ) ? ( in_stream_buff_0 ) : ( in_stream_buff_1 ) ;
assign n305 =  ( n32 ) ? ( in_stream_buff_1 ) : ( n304 ) ;
assign n306 =  ( n25 ) ? ( in_stream_buff_1 ) : ( n305 ) ;
assign n307 =  ( n18 ) ? ( in_stream_buff_1 ) : ( n306 ) ;
assign n308 =  ( n9 ) ? ( in_stream_buff_1 ) : ( n307 ) ;
assign n309 =  ( n4 ) ? ( in_stream_buff_1 ) : ( n308 ) ;
assign n310 =  ( in_stream_full ) == ( 1'd1 )  ;
assign n311 =  ( n310 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n312 =  ( n37 ) ? ( 1'd0 ) : ( in_stream_empty ) ;
assign n313 =  ( n32 ) ? ( n311 ) : ( n312 ) ;
assign n314 =  ( n25 ) ? ( in_stream_empty ) : ( n313 ) ;
assign n315 =  ( n18 ) ? ( in_stream_empty ) : ( n314 ) ;
assign n316 =  ( n9 ) ? ( in_stream_empty ) : ( n315 ) ;
assign n317 =  ( n4 ) ? ( in_stream_empty ) : ( n316 ) ;
assign n318 =  ( in_stream_empty ) == ( 1'd1 )  ;
assign n319 =  ( n318 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n320 =  ( n37 ) ? ( n319 ) : ( in_stream_full ) ;
assign n321 =  ( n32 ) ? ( 1'd0 ) : ( n320 ) ;
assign n322 =  ( n25 ) ? ( in_stream_full ) : ( n321 ) ;
assign n323 =  ( n18 ) ? ( in_stream_full ) : ( n322 ) ;
assign n324 =  ( n9 ) ? ( in_stream_full ) : ( n323 ) ;
assign n325 =  ( n4 ) ? ( in_stream_full ) : ( n324 ) ;
assign n326 =  ( n310 ) ? ( in_stream_buff_1 ) : ( in_stream_buff_0 ) ;
assign n327 =  ( LB2D_proc_w ) == ( 64'd0 )  ;
assign n328 =  (  LB2D_proc_7 [ LB2D_proc_x ] )  ;
assign n329 =  ( LB2D_proc_w ) == ( 64'd1 )  ;
assign n330 =  (  LB2D_proc_0 [ LB2D_proc_x ] )  ;
assign n331 =  ( LB2D_proc_w ) == ( 64'd2 )  ;
assign n332 =  (  LB2D_proc_1 [ LB2D_proc_x ] )  ;
assign n333 =  ( LB2D_proc_w ) == ( 64'd3 )  ;
assign n334 =  (  LB2D_proc_2 [ LB2D_proc_x ] )  ;
assign n335 =  ( LB2D_proc_w ) == ( 64'd4 )  ;
assign n336 =  (  LB2D_proc_3 [ LB2D_proc_x ] )  ;
assign n337 =  ( LB2D_proc_w ) == ( 64'd5 )  ;
assign n338 =  (  LB2D_proc_4 [ LB2D_proc_x ] )  ;
assign n339 =  ( LB2D_proc_w ) == ( 64'd6 )  ;
assign n340 =  (  LB2D_proc_5 [ LB2D_proc_x ] )  ;
assign n341 =  (  LB2D_proc_6 [ LB2D_proc_x ] )  ;
assign n342 =  ( n339 ) ? ( n340 ) : ( n341 ) ;
assign n343 =  ( n337 ) ? ( n338 ) : ( n342 ) ;
assign n344 =  ( n335 ) ? ( n336 ) : ( n343 ) ;
assign n345 =  ( n333 ) ? ( n334 ) : ( n344 ) ;
assign n346 =  ( n331 ) ? ( n332 ) : ( n345 ) ;
assign n347 =  ( n329 ) ? ( n330 ) : ( n346 ) ;
assign n348 =  ( n327 ) ? ( n328 ) : ( n347 ) ;
assign n349 =  ( n339 ) ? ( n338 ) : ( n340 ) ;
assign n350 =  ( n337 ) ? ( n336 ) : ( n349 ) ;
assign n351 =  ( n335 ) ? ( n334 ) : ( n350 ) ;
assign n352 =  ( n333 ) ? ( n332 ) : ( n351 ) ;
assign n353 =  ( n331 ) ? ( n330 ) : ( n352 ) ;
assign n354 =  ( n329 ) ? ( n328 ) : ( n353 ) ;
assign n355 =  ( n327 ) ? ( n341 ) : ( n354 ) ;
assign n356 =  ( n339 ) ? ( n336 ) : ( n338 ) ;
assign n357 =  ( n337 ) ? ( n334 ) : ( n356 ) ;
assign n358 =  ( n335 ) ? ( n332 ) : ( n357 ) ;
assign n359 =  ( n333 ) ? ( n330 ) : ( n358 ) ;
assign n360 =  ( n331 ) ? ( n328 ) : ( n359 ) ;
assign n361 =  ( n329 ) ? ( n341 ) : ( n360 ) ;
assign n362 =  ( n327 ) ? ( n340 ) : ( n361 ) ;
assign n363 =  ( n339 ) ? ( n334 ) : ( n336 ) ;
assign n364 =  ( n337 ) ? ( n332 ) : ( n363 ) ;
assign n365 =  ( n335 ) ? ( n330 ) : ( n364 ) ;
assign n366 =  ( n333 ) ? ( n328 ) : ( n365 ) ;
assign n367 =  ( n331 ) ? ( n341 ) : ( n366 ) ;
assign n368 =  ( n329 ) ? ( n340 ) : ( n367 ) ;
assign n369 =  ( n327 ) ? ( n338 ) : ( n368 ) ;
assign n370 =  ( n339 ) ? ( n332 ) : ( n334 ) ;
assign n371 =  ( n337 ) ? ( n330 ) : ( n370 ) ;
assign n372 =  ( n335 ) ? ( n328 ) : ( n371 ) ;
assign n373 =  ( n333 ) ? ( n341 ) : ( n372 ) ;
assign n374 =  ( n331 ) ? ( n340 ) : ( n373 ) ;
assign n375 =  ( n329 ) ? ( n338 ) : ( n374 ) ;
assign n376 =  ( n327 ) ? ( n336 ) : ( n375 ) ;
assign n377 =  ( n339 ) ? ( n330 ) : ( n332 ) ;
assign n378 =  ( n337 ) ? ( n328 ) : ( n377 ) ;
assign n379 =  ( n335 ) ? ( n341 ) : ( n378 ) ;
assign n380 =  ( n333 ) ? ( n340 ) : ( n379 ) ;
assign n381 =  ( n331 ) ? ( n338 ) : ( n380 ) ;
assign n382 =  ( n329 ) ? ( n336 ) : ( n381 ) ;
assign n383 =  ( n327 ) ? ( n334 ) : ( n382 ) ;
assign n384 =  ( n339 ) ? ( n328 ) : ( n330 ) ;
assign n385 =  ( n337 ) ? ( n341 ) : ( n384 ) ;
assign n386 =  ( n335 ) ? ( n340 ) : ( n385 ) ;
assign n387 =  ( n333 ) ? ( n338 ) : ( n386 ) ;
assign n388 =  ( n331 ) ? ( n336 ) : ( n387 ) ;
assign n389 =  ( n329 ) ? ( n334 ) : ( n388 ) ;
assign n390 =  ( n327 ) ? ( n332 ) : ( n389 ) ;
assign n391 =  ( n339 ) ? ( n341 ) : ( n328 ) ;
assign n392 =  ( n337 ) ? ( n340 ) : ( n391 ) ;
assign n393 =  ( n335 ) ? ( n338 ) : ( n392 ) ;
assign n394 =  ( n333 ) ? ( n336 ) : ( n393 ) ;
assign n395 =  ( n331 ) ? ( n334 ) : ( n394 ) ;
assign n396 =  ( n329 ) ? ( n332 ) : ( n395 ) ;
assign n397 =  ( n327 ) ? ( n330 ) : ( n396 ) ;
assign n398 =  { ( n390 ) , ( n397 ) }  ;
assign n399 =  { ( n383 ) , ( n398 ) }  ;
assign n400 =  { ( n376 ) , ( n399 ) }  ;
assign n401 =  { ( n369 ) , ( n400 ) }  ;
assign n402 =  { ( n362 ) , ( n401 ) }  ;
assign n403 =  { ( n355 ) , ( n402 ) }  ;
assign n404 =  { ( n348 ) , ( n403 ) }  ;
assign n405 =  { ( n326 ) , ( n404 ) }  ;
assign n406 =  ( n30 ) ? ( slice_stream_buff_0 ) : ( n405 ) ;
assign n407 =  ( n37 ) ? ( slice_stream_buff_0 ) : ( slice_stream_buff_0 ) ;
assign n408 =  ( n32 ) ? ( n406 ) : ( n407 ) ;
assign n409 =  ( n25 ) ? ( slice_stream_buff_0 ) : ( n408 ) ;
assign n410 =  ( n18 ) ? ( slice_stream_buff_0 ) : ( n409 ) ;
assign n411 =  ( n9 ) ? ( slice_stream_buff_0 ) : ( n410 ) ;
assign n412 =  ( n4 ) ? ( slice_stream_buff_0 ) : ( n411 ) ;
assign n413 =  ( n30 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n414 =  ( n37 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_1 ) ;
assign n415 =  ( n32 ) ? ( n413 ) : ( n414 ) ;
assign n416 =  ( n25 ) ? ( slice_stream_buff_1 ) : ( n415 ) ;
assign n417 =  ( n18 ) ? ( slice_stream_buff_1 ) : ( n416 ) ;
assign n418 =  ( n9 ) ? ( slice_stream_buff_1 ) : ( n417 ) ;
assign n419 =  ( n4 ) ? ( slice_stream_buff_1 ) : ( n418 ) ;
assign n420 =  ( n93 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n421 =  ( n30 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n422 =  ( n37 ) ? ( slice_stream_empty ) : ( slice_stream_empty ) ;
assign n423 =  ( n32 ) ? ( n421 ) : ( n422 ) ;
assign n424 =  ( n25 ) ? ( n420 ) : ( n423 ) ;
assign n425 =  ( n18 ) ? ( slice_stream_empty ) : ( n424 ) ;
assign n426 =  ( n9 ) ? ( slice_stream_empty ) : ( n425 ) ;
assign n427 =  ( n4 ) ? ( slice_stream_empty ) : ( n426 ) ;
assign n428 =  ( slice_stream_empty ) == ( 1'd1 )  ;
assign n429 =  ( n428 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n430 =  ( n30 ) ? ( 1'd0 ) : ( n429 ) ;
assign n431 =  ( n37 ) ? ( slice_stream_full ) : ( slice_stream_full ) ;
assign n432 =  ( n32 ) ? ( n430 ) : ( n431 ) ;
assign n433 =  ( n25 ) ? ( 1'd0 ) : ( n432 ) ;
assign n434 =  ( n18 ) ? ( slice_stream_full ) : ( n433 ) ;
assign n435 =  ( n9 ) ? ( slice_stream_full ) : ( n434 ) ;
assign n436 =  ( n4 ) ? ( slice_stream_full ) : ( n435 ) ;
assign n437 =  ( LB2D_shift_x ) >= ( 9'd8 )  ;
assign n438 = n94[71:64] ;
assign n439 = LB2D_shift_0[71:64] ;
assign n440 = LB2D_shift_1[71:64] ;
assign n441 = LB2D_shift_2[71:64] ;
assign n442 = LB2D_shift_3[71:64] ;
assign n443 = LB2D_shift_4[71:64] ;
assign n444 = LB2D_shift_5[71:64] ;
assign n445 = LB2D_shift_6[71:64] ;
assign n446 = LB2D_shift_7[71:64] ;
assign n447 =  { ( n445 ) , ( n446 ) }  ;
assign n448 =  { ( n444 ) , ( n447 ) }  ;
assign n449 =  { ( n443 ) , ( n448 ) }  ;
assign n450 =  { ( n442 ) , ( n449 ) }  ;
assign n451 =  { ( n441 ) , ( n450 ) }  ;
assign n452 =  { ( n440 ) , ( n451 ) }  ;
assign n453 =  { ( n439 ) , ( n452 ) }  ;
assign n454 =  { ( n438 ) , ( n453 ) }  ;
assign n455 = n94[63:56] ;
assign n456 = LB2D_shift_0[63:56] ;
assign n457 = LB2D_shift_1[63:56] ;
assign n458 = LB2D_shift_2[63:56] ;
assign n459 = LB2D_shift_3[63:56] ;
assign n460 = LB2D_shift_4[63:56] ;
assign n461 = LB2D_shift_5[63:56] ;
assign n462 = LB2D_shift_6[63:56] ;
assign n463 = LB2D_shift_7[63:56] ;
assign n464 =  { ( n462 ) , ( n463 ) }  ;
assign n465 =  { ( n461 ) , ( n464 ) }  ;
assign n466 =  { ( n460 ) , ( n465 ) }  ;
assign n467 =  { ( n459 ) , ( n466 ) }  ;
assign n468 =  { ( n458 ) , ( n467 ) }  ;
assign n469 =  { ( n457 ) , ( n468 ) }  ;
assign n470 =  { ( n456 ) , ( n469 ) }  ;
assign n471 =  { ( n455 ) , ( n470 ) }  ;
assign n472 = n94[55:48] ;
assign n473 = LB2D_shift_0[55:48] ;
assign n474 = LB2D_shift_1[55:48] ;
assign n475 = LB2D_shift_2[55:48] ;
assign n476 = LB2D_shift_3[55:48] ;
assign n477 = LB2D_shift_4[55:48] ;
assign n478 = LB2D_shift_5[55:48] ;
assign n479 = LB2D_shift_6[55:48] ;
assign n480 = LB2D_shift_7[55:48] ;
assign n481 =  { ( n479 ) , ( n480 ) }  ;
assign n482 =  { ( n478 ) , ( n481 ) }  ;
assign n483 =  { ( n477 ) , ( n482 ) }  ;
assign n484 =  { ( n476 ) , ( n483 ) }  ;
assign n485 =  { ( n475 ) , ( n484 ) }  ;
assign n486 =  { ( n474 ) , ( n485 ) }  ;
assign n487 =  { ( n473 ) , ( n486 ) }  ;
assign n488 =  { ( n472 ) , ( n487 ) }  ;
assign n489 = n94[47:40] ;
assign n490 = LB2D_shift_0[47:40] ;
assign n491 = LB2D_shift_1[47:40] ;
assign n492 = LB2D_shift_2[47:40] ;
assign n493 = LB2D_shift_3[47:40] ;
assign n494 = LB2D_shift_4[47:40] ;
assign n495 = LB2D_shift_5[47:40] ;
assign n496 = LB2D_shift_6[47:40] ;
assign n497 = LB2D_shift_7[47:40] ;
assign n498 =  { ( n496 ) , ( n497 ) }  ;
assign n499 =  { ( n495 ) , ( n498 ) }  ;
assign n500 =  { ( n494 ) , ( n499 ) }  ;
assign n501 =  { ( n493 ) , ( n500 ) }  ;
assign n502 =  { ( n492 ) , ( n501 ) }  ;
assign n503 =  { ( n491 ) , ( n502 ) }  ;
assign n504 =  { ( n490 ) , ( n503 ) }  ;
assign n505 =  { ( n489 ) , ( n504 ) }  ;
assign n506 = n94[39:32] ;
assign n507 = LB2D_shift_0[39:32] ;
assign n508 = LB2D_shift_1[39:32] ;
assign n509 = LB2D_shift_2[39:32] ;
assign n510 = LB2D_shift_3[39:32] ;
assign n511 = LB2D_shift_4[39:32] ;
assign n512 = LB2D_shift_5[39:32] ;
assign n513 = LB2D_shift_6[39:32] ;
assign n514 = LB2D_shift_7[39:32] ;
assign n515 =  { ( n513 ) , ( n514 ) }  ;
assign n516 =  { ( n512 ) , ( n515 ) }  ;
assign n517 =  { ( n511 ) , ( n516 ) }  ;
assign n518 =  { ( n510 ) , ( n517 ) }  ;
assign n519 =  { ( n509 ) , ( n518 ) }  ;
assign n520 =  { ( n508 ) , ( n519 ) }  ;
assign n521 =  { ( n507 ) , ( n520 ) }  ;
assign n522 =  { ( n506 ) , ( n521 ) }  ;
assign n523 = n94[31:24] ;
assign n524 = LB2D_shift_0[31:24] ;
assign n525 = LB2D_shift_1[31:24] ;
assign n526 = LB2D_shift_2[31:24] ;
assign n527 = LB2D_shift_3[31:24] ;
assign n528 = LB2D_shift_4[31:24] ;
assign n529 = LB2D_shift_5[31:24] ;
assign n530 = LB2D_shift_6[31:24] ;
assign n531 = LB2D_shift_7[31:24] ;
assign n532 =  { ( n530 ) , ( n531 ) }  ;
assign n533 =  { ( n529 ) , ( n532 ) }  ;
assign n534 =  { ( n528 ) , ( n533 ) }  ;
assign n535 =  { ( n527 ) , ( n534 ) }  ;
assign n536 =  { ( n526 ) , ( n535 ) }  ;
assign n537 =  { ( n525 ) , ( n536 ) }  ;
assign n538 =  { ( n524 ) , ( n537 ) }  ;
assign n539 =  { ( n523 ) , ( n538 ) }  ;
assign n540 = n94[23:16] ;
assign n541 = LB2D_shift_0[23:16] ;
assign n542 = LB2D_shift_1[23:16] ;
assign n543 = LB2D_shift_2[23:16] ;
assign n544 = LB2D_shift_3[23:16] ;
assign n545 = LB2D_shift_4[23:16] ;
assign n546 = LB2D_shift_5[23:16] ;
assign n547 = LB2D_shift_6[23:16] ;
assign n548 = LB2D_shift_7[23:16] ;
assign n549 =  { ( n547 ) , ( n548 ) }  ;
assign n550 =  { ( n546 ) , ( n549 ) }  ;
assign n551 =  { ( n545 ) , ( n550 ) }  ;
assign n552 =  { ( n544 ) , ( n551 ) }  ;
assign n553 =  { ( n543 ) , ( n552 ) }  ;
assign n554 =  { ( n542 ) , ( n553 ) }  ;
assign n555 =  { ( n541 ) , ( n554 ) }  ;
assign n556 =  { ( n540 ) , ( n555 ) }  ;
assign n557 = n94[15:8] ;
assign n558 = LB2D_shift_0[15:8] ;
assign n559 = LB2D_shift_1[15:8] ;
assign n560 = LB2D_shift_2[15:8] ;
assign n561 = LB2D_shift_3[15:8] ;
assign n562 = LB2D_shift_4[15:8] ;
assign n563 = LB2D_shift_5[15:8] ;
assign n564 = LB2D_shift_6[15:8] ;
assign n565 = LB2D_shift_7[15:8] ;
assign n566 =  { ( n564 ) , ( n565 ) }  ;
assign n567 =  { ( n563 ) , ( n566 ) }  ;
assign n568 =  { ( n562 ) , ( n567 ) }  ;
assign n569 =  { ( n561 ) , ( n568 ) }  ;
assign n570 =  { ( n560 ) , ( n569 ) }  ;
assign n571 =  { ( n559 ) , ( n570 ) }  ;
assign n572 =  { ( n558 ) , ( n571 ) }  ;
assign n573 =  { ( n557 ) , ( n572 ) }  ;
assign n574 = n94[7:0] ;
assign n575 = LB2D_shift_0[7:0] ;
assign n576 = LB2D_shift_1[7:0] ;
assign n577 = LB2D_shift_2[7:0] ;
assign n578 = LB2D_shift_3[7:0] ;
assign n579 = LB2D_shift_4[7:0] ;
assign n580 = LB2D_shift_5[7:0] ;
assign n581 = LB2D_shift_6[7:0] ;
assign n582 = LB2D_shift_7[7:0] ;
assign n583 =  { ( n581 ) , ( n582 ) }  ;
assign n584 =  { ( n580 ) , ( n583 ) }  ;
assign n585 =  { ( n579 ) , ( n584 ) }  ;
assign n586 =  { ( n578 ) , ( n585 ) }  ;
assign n587 =  { ( n577 ) , ( n586 ) }  ;
assign n588 =  { ( n576 ) , ( n587 ) }  ;
assign n589 =  { ( n575 ) , ( n588 ) }  ;
assign n590 =  { ( n574 ) , ( n589 ) }  ;
assign n591 =  { ( n573 ) , ( n590 ) }  ;
assign n592 =  { ( n556 ) , ( n591 ) }  ;
assign n593 =  { ( n539 ) , ( n592 ) }  ;
assign n594 =  { ( n522 ) , ( n593 ) }  ;
assign n595 =  { ( n505 ) , ( n594 ) }  ;
assign n596 =  { ( n488 ) , ( n595 ) }  ;
assign n597 =  { ( n471 ) , ( n596 ) }  ;
assign n598 =  { ( n454 ) , ( n597 ) }  ;
assign n599 =  ( n437 ) ? ( n598 ) : ( stencil_stream_buff_0 ) ;
assign n600 =  ( n37 ) ? ( stencil_stream_buff_0 ) : ( stencil_stream_buff_0 ) ;
assign n601 =  ( n32 ) ? ( stencil_stream_buff_0 ) : ( n600 ) ;
assign n602 =  ( n25 ) ? ( n599 ) : ( n601 ) ;
assign n603 =  ( n18 ) ? ( stencil_stream_buff_0 ) : ( n602 ) ;
assign n604 =  ( n9 ) ? ( stencil_stream_buff_0 ) : ( n603 ) ;
assign n605 =  ( n4 ) ? ( stencil_stream_buff_0 ) : ( n604 ) ;
assign n606 =  ( n37 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_1 ) ;
assign n607 =  ( n32 ) ? ( stencil_stream_buff_1 ) : ( n606 ) ;
assign n608 =  ( n25 ) ? ( stencil_stream_buff_0 ) : ( n607 ) ;
assign n609 =  ( n18 ) ? ( stencil_stream_buff_1 ) : ( n608 ) ;
assign n610 =  ( n9 ) ? ( stencil_stream_buff_1 ) : ( n609 ) ;
assign n611 =  ( n4 ) ? ( stencil_stream_buff_1 ) : ( n610 ) ;
assign n612 =  ( n161 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n613 =  ( n23 ) ? ( stencil_stream_empty ) : ( 1'd0 ) ;
assign n614 =  ( n37 ) ? ( stencil_stream_empty ) : ( stencil_stream_empty ) ;
assign n615 =  ( n32 ) ? ( stencil_stream_empty ) : ( n614 ) ;
assign n616 =  ( n25 ) ? ( n613 ) : ( n615 ) ;
assign n617 =  ( n18 ) ? ( n612 ) : ( n616 ) ;
assign n618 =  ( n9 ) ? ( stencil_stream_empty ) : ( n617 ) ;
assign n619 =  ( n4 ) ? ( stencil_stream_empty ) : ( n618 ) ;
assign n620 =  ( n14 ) ? ( 1'd0 ) : ( 1'd0 ) ;
assign n621 =  ( stencil_stream_empty ) == ( 1'd1 )  ;
assign n622 =  ( n621 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n623 =  ( n23 ) ? ( stencil_stream_full ) : ( n622 ) ;
assign n624 =  ( n37 ) ? ( stencil_stream_full ) : ( stencil_stream_full ) ;
assign n625 =  ( n32 ) ? ( stencil_stream_full ) : ( n624 ) ;
assign n626 =  ( n25 ) ? ( n623 ) : ( n625 ) ;
assign n627 =  ( n18 ) ? ( n620 ) : ( n626 ) ;
assign n628 =  ( n9 ) ? ( stencil_stream_full ) : ( n627 ) ;
assign n629 =  ( n4 ) ? ( stencil_stream_full ) : ( n628 ) ;
assign n630 = ~ ( n4 ) ;
assign n631 = ~ ( n9 ) ;
assign n632 =  ( n630 ) & ( n631 )  ;
assign n633 = ~ ( n18 ) ;
assign n634 =  ( n632 ) & ( n633 )  ;
assign n635 = ~ ( n25 ) ;
assign n636 =  ( n634 ) & ( n635 )  ;
assign n637 = ~ ( n32 ) ;
assign n638 =  ( n636 ) & ( n637 )  ;
assign n639 = ~ ( n37 ) ;
assign n640 =  ( n638 ) & ( n639 )  ;
assign n641 =  ( n638 ) & ( n37 )  ;
assign n642 =  ( n636 ) & ( n32 )  ;
assign n643 = ~ ( n327 ) ;
assign n644 =  ( n642 ) & ( n643 )  ;
assign n645 =  ( n642 ) & ( n327 )  ;
assign n646 =  ( n634 ) & ( n25 )  ;
assign n647 =  ( n632 ) & ( n18 )  ;
assign n648 =  ( n630 ) & ( n9 )  ;
assign LB2D_proc_0_addr0 = n645 ? (LB2D_proc_x) : (0);
assign LB2D_proc_0_data0 = n645 ? (n326) : (LB2D_proc_0[0]);
assign n649 = ~ ( n329 ) ;
assign n650 =  ( n642 ) & ( n649 )  ;
assign n651 =  ( n642 ) & ( n329 )  ;
assign LB2D_proc_1_addr0 = n651 ? (LB2D_proc_x) : (0);
assign LB2D_proc_1_data0 = n651 ? (n326) : (LB2D_proc_1[0]);
assign n652 = ~ ( n331 ) ;
assign n653 =  ( n642 ) & ( n652 )  ;
assign n654 =  ( n642 ) & ( n331 )  ;
assign LB2D_proc_2_addr0 = n654 ? (LB2D_proc_x) : (0);
assign LB2D_proc_2_data0 = n654 ? (n326) : (LB2D_proc_2[0]);
assign n655 = ~ ( n333 ) ;
assign n656 =  ( n642 ) & ( n655 )  ;
assign n657 =  ( n642 ) & ( n333 )  ;
assign LB2D_proc_3_addr0 = n657 ? (LB2D_proc_x) : (0);
assign LB2D_proc_3_data0 = n657 ? (n326) : (LB2D_proc_3[0]);
assign n658 = ~ ( n335 ) ;
assign n659 =  ( n642 ) & ( n658 )  ;
assign n660 =  ( n642 ) & ( n335 )  ;
assign LB2D_proc_4_addr0 = n660 ? (LB2D_proc_x) : (0);
assign LB2D_proc_4_data0 = n660 ? (n326) : (LB2D_proc_4[0]);
assign n661 = ~ ( n337 ) ;
assign n662 =  ( n642 ) & ( n661 )  ;
assign n663 =  ( n642 ) & ( n337 )  ;
assign LB2D_proc_5_addr0 = n663 ? (LB2D_proc_x) : (0);
assign LB2D_proc_5_data0 = n663 ? (n326) : (LB2D_proc_5[0]);
assign n664 = ~ ( n339 ) ;
assign n665 =  ( n642 ) & ( n664 )  ;
assign n666 =  ( n642 ) & ( n339 )  ;
assign LB2D_proc_6_addr0 = n666 ? (LB2D_proc_x) : (0);
assign LB2D_proc_6_data0 = n666 ? (n326) : (LB2D_proc_6[0]);
assign n667 =  ( LB2D_proc_w ) == ( 64'd7 )  ;
assign n668 = ~ ( n667 ) ;
assign n669 =  ( n642 ) & ( n668 )  ;
assign n670 =  ( n642 ) & ( n667 )  ;
assign LB2D_proc_7_addr0 = n670 ? (LB2D_proc_x) : (0);
assign LB2D_proc_7_data0 = n670 ? (n326) : (LB2D_proc_7[0]);
function [7:0] gb_fun ;
input [647:0] arg0;
    begin
//TODO: Add the specific function HERE.    end
endfunction

always @(posedge clk) begin
   if(rst) begin
       LB1D_buff <= LB1D_buff;
       LB1D_in <= LB1D_in;
       LB1D_it_1 <= LB1D_it_1;
       LB1D_p_cnt <= LB1D_p_cnt;
       LB2D_proc_w <= LB2D_proc_w;
       LB2D_proc_x <= LB2D_proc_x;
       LB2D_proc_y <= LB2D_proc_y;
       LB2D_shift_0 <= LB2D_shift_0;
       LB2D_shift_1 <= LB2D_shift_1;
       LB2D_shift_2 <= LB2D_shift_2;
       LB2D_shift_3 <= LB2D_shift_3;
       LB2D_shift_4 <= LB2D_shift_4;
       LB2D_shift_5 <= LB2D_shift_5;
       LB2D_shift_6 <= LB2D_shift_6;
       LB2D_shift_7 <= LB2D_shift_7;
       LB2D_shift_x <= LB2D_shift_x;
       LB2D_shift_y <= LB2D_shift_y;
       arg_0_TDATA <= arg_0_TDATA;
       arg_0_TVALID <= arg_0_TVALID;
       arg_1_TREADY <= arg_1_TREADY;
       gb_exit_it_1 <= gb_exit_it_1;
       gb_exit_it_2 <= gb_exit_it_2;
       gb_exit_it_3 <= gb_exit_it_3;
       gb_exit_it_4 <= gb_exit_it_4;
       gb_exit_it_5 <= gb_exit_it_5;
       gb_exit_it_6 <= gb_exit_it_6;
       gb_exit_it_7 <= gb_exit_it_7;
       gb_exit_it_8 <= gb_exit_it_8;
       gb_p_cnt <= gb_p_cnt;
       gb_pp_it_1 <= gb_pp_it_1;
       gb_pp_it_2 <= gb_pp_it_2;
       gb_pp_it_3 <= gb_pp_it_3;
       gb_pp_it_4 <= gb_pp_it_4;
       gb_pp_it_5 <= gb_pp_it_5;
       gb_pp_it_6 <= gb_pp_it_6;
       gb_pp_it_7 <= gb_pp_it_7;
       gb_pp_it_8 <= gb_pp_it_8;
       gb_pp_it_9 <= gb_pp_it_9;
       in_stream_buff_0 <= in_stream_buff_0;
       in_stream_buff_1 <= in_stream_buff_1;
       in_stream_empty <= in_stream_empty;
       in_stream_full <= in_stream_full;
       slice_stream_buff_0 <= slice_stream_buff_0;
       slice_stream_buff_1 <= slice_stream_buff_1;
       slice_stream_empty <= slice_stream_empty;
       slice_stream_full <= slice_stream_full;
       stencil_stream_buff_0 <= stencil_stream_buff_0;
       stencil_stream_buff_1 <= stencil_stream_buff_1;
       stencil_stream_empty <= stencil_stream_empty;
       stencil_stream_full <= stencil_stream_full;
   end
   else if(step) begin
       LB1D_buff <= n43;
       LB1D_in <= n48;
       LB1D_it_1 <= n51;
       LB1D_p_cnt <= n62;
       LB2D_proc_w <= n73;
       LB2D_proc_x <= n84;
       LB2D_proc_y <= n92;
       LB2D_shift_0 <= n100;
       LB2D_shift_1 <= n106;
       LB2D_shift_2 <= n112;
       LB2D_shift_3 <= n118;
       LB2D_shift_4 <= n124;
       LB2D_shift_5 <= n130;
       LB2D_shift_6 <= n136;
       LB2D_shift_7 <= n142;
       LB2D_shift_x <= n149;
       LB2D_shift_y <= n160;
       arg_0_TDATA <= n169;
       arg_0_TVALID <= n177;
       arg_1_TREADY <= n184;
       gb_exit_it_1 <= n193;
       gb_exit_it_2 <= n199;
       gb_exit_it_3 <= n205;
       gb_exit_it_4 <= n211;
       gb_exit_it_5 <= n217;
       gb_exit_it_6 <= n223;
       gb_exit_it_7 <= n229;
       gb_exit_it_8 <= n235;
       gb_p_cnt <= n243;
       gb_pp_it_1 <= n249;
       gb_pp_it_2 <= n255;
       gb_pp_it_3 <= n261;
       gb_pp_it_4 <= n267;
       gb_pp_it_5 <= n273;
       gb_pp_it_6 <= n279;
       gb_pp_it_7 <= n285;
       gb_pp_it_8 <= n291;
       gb_pp_it_9 <= n297;
       in_stream_buff_0 <= n303;
       in_stream_buff_1 <= n309;
       in_stream_empty <= n317;
       in_stream_full <= n325;
       slice_stream_buff_0 <= n412;
       slice_stream_buff_1 <= n419;
       slice_stream_empty <= n427;
       slice_stream_full <= n436;
       stencil_stream_buff_0 <= n605;
       stencil_stream_buff_1 <= n611;
       stencil_stream_empty <= n619;
       stencil_stream_full <= n629;
       LB2D_proc_0 [ LB2D_proc_0_addr0 ] <= LB2D_proc_0_data0;
       LB2D_proc_1 [ LB2D_proc_1_addr0 ] <= LB2D_proc_1_data0;
       LB2D_proc_2 [ LB2D_proc_2_addr0 ] <= LB2D_proc_2_data0;
       LB2D_proc_3 [ LB2D_proc_3_addr0 ] <= LB2D_proc_3_data0;
       LB2D_proc_4 [ LB2D_proc_4_addr0 ] <= LB2D_proc_4_data0;
       LB2D_proc_5 [ LB2D_proc_5_addr0 ] <= LB2D_proc_5_data0;
       LB2D_proc_6 [ LB2D_proc_6_addr0 ] <= LB2D_proc_6_data0;
       LB2D_proc_7 [ LB2D_proc_7_addr0 ] <= LB2D_proc_7_data0;
   end
end
endmodule
