module GB(
arg_0_TREADY,
arg_1_TDATA,
arg_1_TVALID,
LB1D_buff,
LB1D_it_1,
LB1D_p_cnt,
LB2D_proc_w,
LB2D_proc_x,
LB2D_proc_y,
LB2D_shift_0,
LB2D_shift_1,
LB2D_shift_2,
LB2D_shift_3,
LB2D_shift_4,
LB2D_shift_5,
LB2D_shift_6,
LB2D_shift_7,
LB2D_shift_x,
LB2D_shift_y,
arg_0_TDATA,
arg_0_TVALID,
arg_1_TREADY,
gb_exit_it_1,
gb_exit_it_2,
gb_exit_it_3,
gb_exit_it_4,
gb_exit_it_5,
gb_exit_it_6,
gb_exit_it_7,
gb_exit_it_8,
gb_p_cnt,
gb_pp_it_1,
gb_pp_it_2,
gb_pp_it_3,
gb_pp_it_4,
gb_pp_it_5,
gb_pp_it_6,
gb_pp_it_7,
gb_pp_it_8,
gb_pp_it_9,
in_stream_buff_0,
in_stream_buff_1,
in_stream_empty,
in_stream_full,
slice_stream_buff_0,
slice_stream_buff_1,
slice_stream_empty,
slice_stream_full,
stencil_stream_buff_0,
stencil_stream_buff_1,
stencil_stream_empty,
stencil_stream_full,
clk,rst,
step
);
input            arg_0_TREADY;
input      [7:0] arg_1_TDATA;
input            arg_1_TVALID;
input clk;
input rst;
input step;
output      [7:0] LB1D_buff;
output            LB1D_it_1;
output     [18:0] LB1D_p_cnt;
output     [63:0] LB2D_proc_w;
output      [8:0] LB2D_proc_x;
output      [9:0] LB2D_proc_y;
output     [71:0] LB2D_shift_0;
output     [71:0] LB2D_shift_1;
output     [71:0] LB2D_shift_2;
output     [71:0] LB2D_shift_3;
output     [71:0] LB2D_shift_4;
output     [71:0] LB2D_shift_5;
output     [71:0] LB2D_shift_6;
output     [71:0] LB2D_shift_7;
output      [8:0] LB2D_shift_x;
output      [9:0] LB2D_shift_y;
output      [7:0] arg_0_TDATA;
output            arg_0_TVALID;
output            arg_1_TREADY;
output            gb_exit_it_1;
output            gb_exit_it_2;
output            gb_exit_it_3;
output            gb_exit_it_4;
output            gb_exit_it_5;
output            gb_exit_it_6;
output            gb_exit_it_7;
output            gb_exit_it_8;
output     [18:0] gb_p_cnt;
output            gb_pp_it_1;
output            gb_pp_it_2;
output            gb_pp_it_3;
output            gb_pp_it_4;
output            gb_pp_it_5;
output            gb_pp_it_6;
output            gb_pp_it_7;
output            gb_pp_it_8;
output            gb_pp_it_9;
output      [7:0] in_stream_buff_0;
output      [7:0] in_stream_buff_1;
output            in_stream_empty;
output            in_stream_full;
output     [71:0] slice_stream_buff_0;
output     [71:0] slice_stream_buff_1;
output            slice_stream_empty;
output            slice_stream_full;
output    [647:0] stencil_stream_buff_0;
output    [647:0] stencil_stream_buff_1;
output            stencil_stream_empty;
output            stencil_stream_full;
reg      [7:0] LB1D_buff;
reg            LB1D_it_1;
reg     [18:0] LB1D_p_cnt;
reg     [63:0] LB2D_proc_w;
reg      [8:0] LB2D_proc_x;
reg      [9:0] LB2D_proc_y;
reg     [71:0] LB2D_shift_0;
reg     [71:0] LB2D_shift_1;
reg     [71:0] LB2D_shift_2;
reg     [71:0] LB2D_shift_3;
reg     [71:0] LB2D_shift_4;
reg     [71:0] LB2D_shift_5;
reg     [71:0] LB2D_shift_6;
reg     [71:0] LB2D_shift_7;
reg      [8:0] LB2D_shift_x;
reg      [9:0] LB2D_shift_y;
reg      [7:0] arg_0_TDATA;
reg            arg_0_TVALID;
reg            arg_1_TREADY;
reg            gb_exit_it_1;
reg            gb_exit_it_2;
reg            gb_exit_it_3;
reg            gb_exit_it_4;
reg            gb_exit_it_5;
reg            gb_exit_it_6;
reg            gb_exit_it_7;
reg            gb_exit_it_8;
reg     [18:0] gb_p_cnt;
reg            gb_pp_it_1;
reg            gb_pp_it_2;
reg            gb_pp_it_3;
reg            gb_pp_it_4;
reg            gb_pp_it_5;
reg            gb_pp_it_6;
reg            gb_pp_it_7;
reg            gb_pp_it_8;
reg            gb_pp_it_9;
reg      [7:0] in_stream_buff_0;
reg      [7:0] in_stream_buff_1;
reg            in_stream_empty;
reg            in_stream_full;
reg     [71:0] slice_stream_buff_0;
reg     [71:0] slice_stream_buff_1;
reg            slice_stream_empty;
reg            slice_stream_full;
reg    [647:0] stencil_stream_buff_0;
reg    [647:0] stencil_stream_buff_1;
reg            stencil_stream_empty;
reg            stencil_stream_full;
wire            arg_0_TREADY;
wire      [7:0] arg_1_TDATA;
wire            arg_1_TVALID;
wire            n0;
wire            n1;
wire            n2;
wire            n3;
wire            n4;
wire            n5;
wire            n6;
wire            n7;
wire            n8;
wire            n9;
wire            n10;
wire            n11;
wire            n12;
wire            n13;
wire            n14;
wire            n15;
wire            n16;
wire            n17;
wire            n18;
wire            n19;
wire            n20;
wire            n21;
wire            n22;
wire            n23;
wire            n24;
wire            n25;
wire            n26;
wire            n27;
wire            n28;
wire            n29;
wire            n30;
wire            n31;
wire            n32;
wire            n33;
wire            n34;
wire            n35;
wire            n36;
wire            n37;
wire            n38;
wire            n39;
wire      [7:0] n40;
wire      [7:0] n41;
wire      [7:0] n42;
wire      [7:0] n43;
wire      [7:0] n44;
wire      [7:0] n45;
wire            n46;
wire            n47;
wire            n48;
wire     [18:0] n49;
wire     [18:0] n50;
wire     [18:0] n51;
wire     [18:0] n52;
wire     [18:0] n53;
wire     [18:0] n54;
wire     [18:0] n55;
wire     [18:0] n56;
wire            n57;
wire            n58;
wire     [63:0] n59;
wire     [63:0] n60;
wire     [63:0] n61;
wire     [63:0] n62;
wire     [63:0] n63;
wire     [63:0] n64;
wire     [63:0] n65;
wire     [63:0] n66;
wire     [63:0] n67;
wire            n68;
wire            n69;
wire            n70;
wire      [8:0] n71;
wire      [8:0] n72;
wire      [8:0] n73;
wire      [8:0] n74;
wire      [8:0] n75;
wire      [8:0] n76;
wire      [8:0] n77;
wire      [8:0] n78;
wire            n79;
wire      [9:0] n80;
wire      [9:0] n81;
wire      [9:0] n82;
wire      [9:0] n83;
wire      [9:0] n84;
wire      [9:0] n85;
wire      [9:0] n86;
wire            n87;
wire     [71:0] n88;
wire     [71:0] n89;
wire     [71:0] n90;
wire     [71:0] n91;
wire     [71:0] n92;
wire     [71:0] n93;
wire     [71:0] n94;
wire     [71:0] n95;
wire     [71:0] n96;
wire     [71:0] n97;
wire     [71:0] n98;
wire     [71:0] n99;
wire     [71:0] n100;
wire     [71:0] n101;
wire     [71:0] n102;
wire     [71:0] n103;
wire     [71:0] n104;
wire     [71:0] n105;
wire     [71:0] n106;
wire     [71:0] n107;
wire     [71:0] n108;
wire     [71:0] n109;
wire     [71:0] n110;
wire     [71:0] n111;
wire     [71:0] n112;
wire     [71:0] n113;
wire     [71:0] n114;
wire     [71:0] n115;
wire     [71:0] n116;
wire     [71:0] n117;
wire     [71:0] n118;
wire     [71:0] n119;
wire     [71:0] n120;
wire     [71:0] n121;
wire     [71:0] n122;
wire     [71:0] n123;
wire     [71:0] n124;
wire     [71:0] n125;
wire     [71:0] n126;
wire     [71:0] n127;
wire     [71:0] n128;
wire     [71:0] n129;
wire     [71:0] n130;
wire     [71:0] n131;
wire     [71:0] n132;
wire     [71:0] n133;
wire     [71:0] n134;
wire     [71:0] n135;
wire     [71:0] n136;
wire      [8:0] n137;
wire      [8:0] n138;
wire      [8:0] n139;
wire      [8:0] n140;
wire      [8:0] n141;
wire      [8:0] n142;
wire      [8:0] n143;
wire            n144;
wire            n145;
wire      [9:0] n146;
wire      [9:0] n147;
wire      [9:0] n148;
wire      [9:0] n149;
wire      [9:0] n150;
wire      [9:0] n151;
wire      [9:0] n152;
wire      [9:0] n153;
wire      [9:0] n154;
wire            n155;
wire    [647:0] n156;
wire      [7:0] n157;
wire      [7:0] n158;
wire      [7:0] n159;
wire      [7:0] n160;
wire      [7:0] n161;
wire      [7:0] n162;
wire      [7:0] n163;
wire            n164;
wire            n165;
wire            n166;
wire            n167;
wire            n168;
wire            n169;
wire            n170;
wire            n171;
wire            n172;
wire            n173;
wire            n174;
wire            n175;
wire            n176;
wire            n177;
wire            n178;
wire     [18:0] n179;
wire            n180;
wire            n181;
wire            n182;
wire            n183;
wire            n184;
wire            n185;
wire            n186;
wire            n187;
wire            n188;
wire            n189;
wire            n190;
wire            n191;
wire            n192;
wire            n193;
wire            n194;
wire            n195;
wire            n196;
wire            n197;
wire            n198;
wire            n199;
wire            n200;
wire            n201;
wire            n202;
wire            n203;
wire            n204;
wire            n205;
wire            n206;
wire            n207;
wire            n208;
wire            n209;
wire            n210;
wire            n211;
wire            n212;
wire            n213;
wire            n214;
wire            n215;
wire            n216;
wire            n217;
wire            n218;
wire            n219;
wire            n220;
wire            n221;
wire            n222;
wire            n223;
wire            n224;
wire            n225;
wire            n226;
wire            n227;
wire            n228;
wire            n229;
wire            n230;
wire     [18:0] n231;
wire     [18:0] n232;
wire     [18:0] n233;
wire     [18:0] n234;
wire     [18:0] n235;
wire     [18:0] n236;
wire     [18:0] n237;
wire            n238;
wire            n239;
wire            n240;
wire            n241;
wire            n242;
wire            n243;
wire            n244;
wire            n245;
wire            n246;
wire            n247;
wire            n248;
wire            n249;
wire            n250;
wire            n251;
wire            n252;
wire            n253;
wire            n254;
wire            n255;
wire            n256;
wire            n257;
wire            n258;
wire            n259;
wire            n260;
wire            n261;
wire            n262;
wire            n263;
wire            n264;
wire            n265;
wire            n266;
wire            n267;
wire            n268;
wire            n269;
wire            n270;
wire            n271;
wire            n272;
wire            n273;
wire            n274;
wire            n275;
wire            n276;
wire            n277;
wire            n278;
wire            n279;
wire            n280;
wire            n281;
wire            n282;
wire            n283;
wire            n284;
wire            n285;
wire            n286;
wire            n287;
wire            n288;
wire            n289;
wire            n290;
wire            n291;
wire      [7:0] n292;
wire      [7:0] n293;
wire      [7:0] n294;
wire      [7:0] n295;
wire      [7:0] n296;
wire      [7:0] n297;
wire      [7:0] n298;
wire      [7:0] n299;
wire      [7:0] n300;
wire      [7:0] n301;
wire      [7:0] n302;
wire      [7:0] n303;
wire            n304;
wire            n305;
wire            n306;
wire            n307;
wire            n308;
wire            n309;
wire            n310;
wire            n311;
wire            n312;
wire            n313;
wire            n314;
wire            n315;
wire            n316;
wire            n317;
wire            n318;
wire            n319;
wire      [7:0] n320;
wire            n321;
wire      [7:0] n322;
wire            n323;
wire      [7:0] n324;
wire            n325;
wire      [7:0] n326;
wire            n327;
wire      [7:0] n328;
wire            n329;
wire      [7:0] n330;
wire            n331;
wire      [7:0] n332;
wire            n333;
wire      [7:0] n334;
wire      [7:0] n335;
wire      [7:0] n336;
wire      [7:0] n337;
wire      [7:0] n338;
wire      [7:0] n339;
wire      [7:0] n340;
wire      [7:0] n341;
wire      [7:0] n342;
wire      [7:0] n343;
wire      [7:0] n344;
wire      [7:0] n345;
wire      [7:0] n346;
wire      [7:0] n347;
wire      [7:0] n348;
wire      [7:0] n349;
wire      [7:0] n350;
wire      [7:0] n351;
wire      [7:0] n352;
wire      [7:0] n353;
wire      [7:0] n354;
wire      [7:0] n355;
wire      [7:0] n356;
wire      [7:0] n357;
wire      [7:0] n358;
wire      [7:0] n359;
wire      [7:0] n360;
wire      [7:0] n361;
wire      [7:0] n362;
wire      [7:0] n363;
wire      [7:0] n364;
wire      [7:0] n365;
wire      [7:0] n366;
wire      [7:0] n367;
wire      [7:0] n368;
wire      [7:0] n369;
wire      [7:0] n370;
wire      [7:0] n371;
wire      [7:0] n372;
wire      [7:0] n373;
wire      [7:0] n374;
wire      [7:0] n375;
wire      [7:0] n376;
wire      [7:0] n377;
wire      [7:0] n378;
wire      [7:0] n379;
wire      [7:0] n380;
wire      [7:0] n381;
wire      [7:0] n382;
wire      [7:0] n383;
wire      [7:0] n384;
wire      [7:0] n385;
wire      [7:0] n386;
wire      [7:0] n387;
wire      [7:0] n388;
wire      [7:0] n389;
wire      [7:0] n390;
wire      [7:0] n391;
wire     [15:0] n392;
wire     [23:0] n393;
wire     [31:0] n394;
wire     [39:0] n395;
wire     [47:0] n396;
wire     [55:0] n397;
wire     [63:0] n398;
wire     [71:0] n399;
wire     [71:0] n400;
wire     [71:0] n401;
wire     [71:0] n402;
wire     [71:0] n403;
wire     [71:0] n404;
wire     [71:0] n405;
wire     [71:0] n406;
wire     [71:0] n407;
wire     [71:0] n408;
wire     [71:0] n409;
wire     [71:0] n410;
wire     [71:0] n411;
wire     [71:0] n412;
wire     [71:0] n413;
wire            n414;
wire            n415;
wire            n416;
wire            n417;
wire            n418;
wire            n419;
wire            n420;
wire            n421;
wire            n422;
wire            n423;
wire            n424;
wire            n425;
wire            n426;
wire            n427;
wire            n428;
wire            n429;
wire            n430;
wire            n431;
wire      [7:0] n432;
wire      [7:0] n433;
wire      [7:0] n434;
wire      [7:0] n435;
wire      [7:0] n436;
wire      [7:0] n437;
wire      [7:0] n438;
wire      [7:0] n439;
wire      [7:0] n440;
wire     [15:0] n441;
wire     [23:0] n442;
wire     [31:0] n443;
wire     [39:0] n444;
wire     [47:0] n445;
wire     [55:0] n446;
wire     [63:0] n447;
wire     [71:0] n448;
wire      [7:0] n449;
wire      [7:0] n450;
wire      [7:0] n451;
wire      [7:0] n452;
wire      [7:0] n453;
wire      [7:0] n454;
wire      [7:0] n455;
wire      [7:0] n456;
wire      [7:0] n457;
wire     [15:0] n458;
wire     [23:0] n459;
wire     [31:0] n460;
wire     [39:0] n461;
wire     [47:0] n462;
wire     [55:0] n463;
wire     [63:0] n464;
wire     [71:0] n465;
wire      [7:0] n466;
wire      [7:0] n467;
wire      [7:0] n468;
wire      [7:0] n469;
wire      [7:0] n470;
wire      [7:0] n471;
wire      [7:0] n472;
wire      [7:0] n473;
wire      [7:0] n474;
wire     [15:0] n475;
wire     [23:0] n476;
wire     [31:0] n477;
wire     [39:0] n478;
wire     [47:0] n479;
wire     [55:0] n480;
wire     [63:0] n481;
wire     [71:0] n482;
wire      [7:0] n483;
wire      [7:0] n484;
wire      [7:0] n485;
wire      [7:0] n486;
wire      [7:0] n487;
wire      [7:0] n488;
wire      [7:0] n489;
wire      [7:0] n490;
wire      [7:0] n491;
wire     [15:0] n492;
wire     [23:0] n493;
wire     [31:0] n494;
wire     [39:0] n495;
wire     [47:0] n496;
wire     [55:0] n497;
wire     [63:0] n498;
wire     [71:0] n499;
wire      [7:0] n500;
wire      [7:0] n501;
wire      [7:0] n502;
wire      [7:0] n503;
wire      [7:0] n504;
wire      [7:0] n505;
wire      [7:0] n506;
wire      [7:0] n507;
wire      [7:0] n508;
wire     [15:0] n509;
wire     [23:0] n510;
wire     [31:0] n511;
wire     [39:0] n512;
wire     [47:0] n513;
wire     [55:0] n514;
wire     [63:0] n515;
wire     [71:0] n516;
wire      [7:0] n517;
wire      [7:0] n518;
wire      [7:0] n519;
wire      [7:0] n520;
wire      [7:0] n521;
wire      [7:0] n522;
wire      [7:0] n523;
wire      [7:0] n524;
wire      [7:0] n525;
wire     [15:0] n526;
wire     [23:0] n527;
wire     [31:0] n528;
wire     [39:0] n529;
wire     [47:0] n530;
wire     [55:0] n531;
wire     [63:0] n532;
wire     [71:0] n533;
wire      [7:0] n534;
wire      [7:0] n535;
wire      [7:0] n536;
wire      [7:0] n537;
wire      [7:0] n538;
wire      [7:0] n539;
wire      [7:0] n540;
wire      [7:0] n541;
wire      [7:0] n542;
wire     [15:0] n543;
wire     [23:0] n544;
wire     [31:0] n545;
wire     [39:0] n546;
wire     [47:0] n547;
wire     [55:0] n548;
wire     [63:0] n549;
wire     [71:0] n550;
wire      [7:0] n551;
wire      [7:0] n552;
wire      [7:0] n553;
wire      [7:0] n554;
wire      [7:0] n555;
wire      [7:0] n556;
wire      [7:0] n557;
wire      [7:0] n558;
wire      [7:0] n559;
wire     [15:0] n560;
wire     [23:0] n561;
wire     [31:0] n562;
wire     [39:0] n563;
wire     [47:0] n564;
wire     [55:0] n565;
wire     [63:0] n566;
wire     [71:0] n567;
wire      [7:0] n568;
wire      [7:0] n569;
wire      [7:0] n570;
wire      [7:0] n571;
wire      [7:0] n572;
wire      [7:0] n573;
wire      [7:0] n574;
wire      [7:0] n575;
wire      [7:0] n576;
wire     [15:0] n577;
wire     [23:0] n578;
wire     [31:0] n579;
wire     [39:0] n580;
wire     [47:0] n581;
wire     [55:0] n582;
wire     [63:0] n583;
wire     [71:0] n584;
wire    [143:0] n585;
wire    [215:0] n586;
wire    [287:0] n587;
wire    [359:0] n588;
wire    [431:0] n589;
wire    [503:0] n590;
wire    [575:0] n591;
wire    [647:0] n592;
wire    [647:0] n593;
wire    [647:0] n594;
wire    [647:0] n595;
wire    [647:0] n596;
wire    [647:0] n597;
wire    [647:0] n598;
wire    [647:0] n599;
wire    [647:0] n600;
wire    [647:0] n601;
wire    [647:0] n602;
wire    [647:0] n603;
wire    [647:0] n604;
wire    [647:0] n605;
wire            n606;
wire            n607;
wire            n608;
wire            n609;
wire            n610;
wire            n611;
wire            n612;
wire            n613;
wire            n614;
wire            n615;
wire            n616;
wire            n617;
wire            n618;
wire            n619;
wire            n620;
wire            n621;
wire            n622;
wire            n623;
wire      [8:0] LB2D_proc_0_addr0;
wire      [7:0] LB2D_proc_0_data0;
wire            n624;
wire            n625;
wire            n626;
wire            n627;
wire            n628;
wire            n629;
wire            n630;
wire            n631;
wire            n632;
wire            n633;
wire            n634;
wire            n635;
wire            n636;
wire            n637;
wire            n638;
wire            n639;
wire            n640;
wire            n641;
wire            n642;
wire      [8:0] LB2D_proc_1_addr0;
wire      [7:0] LB2D_proc_1_data0;
wire            n643;
wire            n644;
wire            n645;
wire      [8:0] LB2D_proc_2_addr0;
wire      [7:0] LB2D_proc_2_data0;
wire            n646;
wire            n647;
wire            n648;
wire      [8:0] LB2D_proc_3_addr0;
wire      [7:0] LB2D_proc_3_data0;
wire            n649;
wire            n650;
wire            n651;
wire      [8:0] LB2D_proc_4_addr0;
wire      [7:0] LB2D_proc_4_data0;
wire            n652;
wire            n653;
wire            n654;
wire      [8:0] LB2D_proc_5_addr0;
wire      [7:0] LB2D_proc_5_data0;
wire            n655;
wire            n656;
wire            n657;
wire      [8:0] LB2D_proc_6_addr0;
wire      [7:0] LB2D_proc_6_data0;
wire            n658;
wire            n659;
wire            n660;
wire      [8:0] LB2D_proc_7_addr0;
wire      [7:0] LB2D_proc_7_data0;
wire            n661;
wire            n662;
wire            n663;
wire            n664;
reg      [7:0] LB2D_proc_0[511:0];
reg      [7:0] LB2D_proc_1[511:0];
reg      [7:0] LB2D_proc_2[511:0];
reg      [7:0] LB2D_proc_3[511:0];
reg      [7:0] LB2D_proc_4[511:0];
reg      [7:0] LB2D_proc_5[511:0];
reg      [7:0] LB2D_proc_6[511:0];
reg      [7:0] LB2D_proc_7[511:0];
wire clk;
wire rst;
wire step;
assign n0 =  ( arg_0_TREADY ) == ( 1'd1 )  ;
assign n1 =  ( arg_0_TVALID ) == ( 1'd1 )  ;
assign n2 =  ( n0 ) & ( n1 )  ;
assign n3 =  ( arg_1_TVALID ) == ( 1'd0 )  ;
assign n4 =  ( n2 ) & ( n3 )  ;
assign n5 =  ( arg_1_TREADY ) == ( 1'd1 )  ;
assign n6 =  ( arg_1_TVALID ) == ( 1'd1 )  ;
assign n7 =  ( n5 ) & ( n6 )  ;
assign n8 =  ( arg_0_TREADY ) == ( 1'd0 )  ;
assign n9 =  ( n7 ) & ( n8 )  ;
assign n10 =  ( arg_0_TVALID ) == ( 1'd0 )  ;
assign n11 =  ( gb_exit_it_1 ) == ( 1'd0 )  ;
assign n12 =  ( stencil_stream_empty ) == ( 1'd0 )  ;
assign n13 =  ( n11 ) & ( n12 )  ;
assign n14 =  ( gb_exit_it_1 ) == ( 1'd1 )  ;
assign n15 =  ( gb_exit_it_8 ) == ( 1'd0 )  ;
assign n16 =  ( n14 ) & ( n15 )  ;
assign n17 =  ( n13 ) | ( n16 )  ;
assign n18 =  ( n10 ) & ( n17 )  ;
assign n19 =  ( slice_stream_empty ) == ( 1'd0 )  ;
assign n20 =  ( LB2D_shift_x ) != ( 9'd488 )  ;
assign n21 =  ( n19 ) & ( n20 )  ;
assign n22 =  ( stencil_stream_full ) == ( 1'd0 )  ;
assign n23 =  ( LB2D_shift_x ) < ( 9'd8 )  ;
assign n24 =  ( n22 ) | ( n23 )  ;
assign n25 =  ( n21 ) & ( n24 )  ;
assign n26 =  ( in_stream_empty ) == ( 1'd0 )  ;
assign n27 =  ( LB2D_proc_x ) != ( 9'd488 )  ;
assign n28 =  ( n26 ) & ( n27 )  ;
assign n29 =  ( slice_stream_full ) == ( 1'd0 )  ;
assign n30 =  ( LB2D_proc_y ) < ( 10'd8 )  ;
assign n31 =  ( n29 ) | ( n30 )  ;
assign n32 =  ( n28 ) & ( n31 )  ;
assign n33 =  ( arg_1_TREADY ) == ( 1'd0 )  ;
assign n34 =  ( in_stream_full ) == ( 1'd0 )  ;
assign n35 =  ( n33 ) & ( n34 )  ;
assign n36 =  ( LB1D_p_cnt ) != ( 19'd316224 )  ;
assign n37 =  ( n35 ) & ( n36 )  ;
assign n38 =  ( LB1D_it_1 ) == ( 1'd1 )  ;
assign n39 =  ( n37 ) & ( n38 )  ;
assign n40 =  ( n39 ) ? ( LB1D_buff ) : ( LB1D_buff ) ;
assign n41 =  ( n32 ) ? ( LB1D_buff ) : ( n40 ) ;
assign n42 =  ( n25 ) ? ( LB1D_buff ) : ( n41 ) ;
assign n43 =  ( n18 ) ? ( LB1D_buff ) : ( n42 ) ;
assign n44 =  ( n9 ) ? ( arg_1_TDATA ) : ( n43 ) ;
assign n45 =  ( n4 ) ? ( arg_1_TDATA ) : ( n44 ) ;
assign n46 =  ( LB1D_it_1 ) == ( 1'd0 )  ;
assign n47 =  ( n37 ) & ( n46 )  ;
assign n48 =  ( n47 ) ? ( 1'd1 ) : ( LB1D_it_1 ) ;
assign n49 =  ( LB1D_p_cnt ) + ( 19'd1 )  ;
assign n50 =  ( n39 ) ? ( n49 ) : ( LB1D_p_cnt ) ;
assign n51 =  ( n47 ) ? ( n49 ) : ( n50 ) ;
assign n52 =  ( n32 ) ? ( LB1D_p_cnt ) : ( n51 ) ;
assign n53 =  ( n25 ) ? ( LB1D_p_cnt ) : ( n52 ) ;
assign n54 =  ( n18 ) ? ( LB1D_p_cnt ) : ( n53 ) ;
assign n55 =  ( n9 ) ? ( LB1D_p_cnt ) : ( n54 ) ;
assign n56 =  ( n4 ) ? ( LB1D_p_cnt ) : ( n55 ) ;
assign n57 =  ( LB2D_proc_w ) < ( 64'd7 )  ;
assign n58 =  ( LB2D_proc_x ) < ( 9'd488 )  ;
assign n59 =  ( LB2D_proc_w ) + ( 64'd1 )  ;
assign n60 =  ( n58 ) ? ( LB2D_proc_w ) : ( n59 ) ;
assign n61 =  ( n57 ) ? ( n60 ) : ( 64'd0 ) ;
assign n62 =  ( n39 ) ? ( LB2D_proc_w ) : ( LB2D_proc_w ) ;
assign n63 =  ( n32 ) ? ( n61 ) : ( n62 ) ;
assign n64 =  ( n25 ) ? ( LB2D_proc_w ) : ( n63 ) ;
assign n65 =  ( n18 ) ? ( LB2D_proc_w ) : ( n64 ) ;
assign n66 =  ( n9 ) ? ( LB2D_proc_w ) : ( n65 ) ;
assign n67 =  ( n4 ) ? ( LB2D_proc_w ) : ( n66 ) ;
assign n68 =  ( LB2D_proc_x ) == ( 9'd488 )  ;
assign n69 =  ( n26 ) & ( n68 )  ;
assign n70 =  ( n69 ) & ( n31 )  ;
assign n71 =  ( LB2D_proc_x ) + ( 9'd1 )  ;
assign n72 =  ( n39 ) ? ( LB2D_proc_x ) : ( LB2D_proc_x ) ;
assign n73 =  ( n32 ) ? ( n71 ) : ( n72 ) ;
assign n74 =  ( n70 ) ? ( 9'd0 ) : ( n73 ) ;
assign n75 =  ( n25 ) ? ( LB2D_proc_x ) : ( n74 ) ;
assign n76 =  ( n18 ) ? ( LB2D_proc_x ) : ( n75 ) ;
assign n77 =  ( n9 ) ? ( LB2D_proc_x ) : ( n76 ) ;
assign n78 =  ( n4 ) ? ( LB2D_proc_x ) : ( n77 ) ;
assign n79 =  ( LB2D_proc_y ) < ( 10'd488 )  ;
assign n80 =  ( n79 ) ? ( LB2D_proc_y ) : ( 10'd488 ) ;
assign n81 =  ( n39 ) ? ( LB2D_proc_y ) : ( LB2D_proc_y ) ;
assign n82 =  ( n32 ) ? ( n80 ) : ( n81 ) ;
assign n83 =  ( n25 ) ? ( LB2D_proc_y ) : ( n82 ) ;
assign n84 =  ( n18 ) ? ( LB2D_proc_y ) : ( n83 ) ;
assign n85 =  ( n9 ) ? ( LB2D_proc_y ) : ( n84 ) ;
assign n86 =  ( n4 ) ? ( LB2D_proc_y ) : ( n85 ) ;
assign n87 =  ( slice_stream_full ) == ( 1'd1 )  ;
assign n88 =  ( n87 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n89 =  ( n39 ) ? ( LB2D_shift_0 ) : ( LB2D_shift_0 ) ;
assign n90 =  ( n32 ) ? ( LB2D_shift_0 ) : ( n89 ) ;
assign n91 =  ( n25 ) ? ( n88 ) : ( n90 ) ;
assign n92 =  ( n18 ) ? ( LB2D_shift_0 ) : ( n91 ) ;
assign n93 =  ( n9 ) ? ( LB2D_shift_0 ) : ( n92 ) ;
assign n94 =  ( n4 ) ? ( LB2D_shift_0 ) : ( n93 ) ;
assign n95 =  ( n39 ) ? ( LB2D_shift_1 ) : ( LB2D_shift_1 ) ;
assign n96 =  ( n32 ) ? ( LB2D_shift_1 ) : ( n95 ) ;
assign n97 =  ( n25 ) ? ( LB2D_shift_0 ) : ( n96 ) ;
assign n98 =  ( n18 ) ? ( LB2D_shift_1 ) : ( n97 ) ;
assign n99 =  ( n9 ) ? ( LB2D_shift_1 ) : ( n98 ) ;
assign n100 =  ( n4 ) ? ( LB2D_shift_1 ) : ( n99 ) ;
assign n101 =  ( n39 ) ? ( LB2D_shift_2 ) : ( LB2D_shift_2 ) ;
assign n102 =  ( n32 ) ? ( LB2D_shift_2 ) : ( n101 ) ;
assign n103 =  ( n25 ) ? ( LB2D_shift_1 ) : ( n102 ) ;
assign n104 =  ( n18 ) ? ( LB2D_shift_2 ) : ( n103 ) ;
assign n105 =  ( n9 ) ? ( LB2D_shift_2 ) : ( n104 ) ;
assign n106 =  ( n4 ) ? ( LB2D_shift_2 ) : ( n105 ) ;
assign n107 =  ( n39 ) ? ( LB2D_shift_3 ) : ( LB2D_shift_3 ) ;
assign n108 =  ( n32 ) ? ( LB2D_shift_3 ) : ( n107 ) ;
assign n109 =  ( n25 ) ? ( LB2D_shift_2 ) : ( n108 ) ;
assign n110 =  ( n18 ) ? ( LB2D_shift_3 ) : ( n109 ) ;
assign n111 =  ( n9 ) ? ( LB2D_shift_3 ) : ( n110 ) ;
assign n112 =  ( n4 ) ? ( LB2D_shift_3 ) : ( n111 ) ;
assign n113 =  ( n39 ) ? ( LB2D_shift_4 ) : ( LB2D_shift_4 ) ;
assign n114 =  ( n32 ) ? ( LB2D_shift_4 ) : ( n113 ) ;
assign n115 =  ( n25 ) ? ( LB2D_shift_3 ) : ( n114 ) ;
assign n116 =  ( n18 ) ? ( LB2D_shift_4 ) : ( n115 ) ;
assign n117 =  ( n9 ) ? ( LB2D_shift_4 ) : ( n116 ) ;
assign n118 =  ( n4 ) ? ( LB2D_shift_4 ) : ( n117 ) ;
assign n119 =  ( n39 ) ? ( LB2D_shift_5 ) : ( LB2D_shift_5 ) ;
assign n120 =  ( n32 ) ? ( LB2D_shift_5 ) : ( n119 ) ;
assign n121 =  ( n25 ) ? ( LB2D_shift_4 ) : ( n120 ) ;
assign n122 =  ( n18 ) ? ( LB2D_shift_5 ) : ( n121 ) ;
assign n123 =  ( n9 ) ? ( LB2D_shift_5 ) : ( n122 ) ;
assign n124 =  ( n4 ) ? ( LB2D_shift_5 ) : ( n123 ) ;
assign n125 =  ( n39 ) ? ( LB2D_shift_6 ) : ( LB2D_shift_6 ) ;
assign n126 =  ( n32 ) ? ( LB2D_shift_6 ) : ( n125 ) ;
assign n127 =  ( n25 ) ? ( LB2D_shift_5 ) : ( n126 ) ;
assign n128 =  ( n18 ) ? ( LB2D_shift_6 ) : ( n127 ) ;
assign n129 =  ( n9 ) ? ( LB2D_shift_6 ) : ( n128 ) ;
assign n130 =  ( n4 ) ? ( LB2D_shift_6 ) : ( n129 ) ;
assign n131 =  ( n39 ) ? ( LB2D_shift_7 ) : ( LB2D_shift_7 ) ;
assign n132 =  ( n32 ) ? ( LB2D_shift_7 ) : ( n131 ) ;
assign n133 =  ( n25 ) ? ( LB2D_shift_6 ) : ( n132 ) ;
assign n134 =  ( n18 ) ? ( LB2D_shift_7 ) : ( n133 ) ;
assign n135 =  ( n9 ) ? ( LB2D_shift_7 ) : ( n134 ) ;
assign n136 =  ( n4 ) ? ( LB2D_shift_7 ) : ( n135 ) ;
assign n137 =  ( LB2D_shift_x ) + ( 9'd1 )  ;
assign n138 =  ( n39 ) ? ( LB2D_shift_x ) : ( LB2D_shift_x ) ;
assign n139 =  ( n32 ) ? ( LB2D_shift_x ) : ( n138 ) ;
assign n140 =  ( n25 ) ? ( n137 ) : ( n139 ) ;
assign n141 =  ( n18 ) ? ( LB2D_shift_x ) : ( n140 ) ;
assign n142 =  ( n9 ) ? ( LB2D_shift_x ) : ( n141 ) ;
assign n143 =  ( n4 ) ? ( LB2D_shift_x ) : ( n142 ) ;
assign n144 =  ( LB2D_shift_y ) < ( 10'd480 )  ;
assign n145 =  ( LB2D_shift_x ) < ( 9'd488 )  ;
assign n146 =  ( LB2D_shift_y ) + ( 10'd1 )  ;
assign n147 =  ( n145 ) ? ( LB2D_shift_y ) : ( n146 ) ;
assign n148 =  ( n144 ) ? ( n147 ) : ( 10'd480 ) ;
assign n149 =  ( n39 ) ? ( LB2D_shift_y ) : ( LB2D_shift_y ) ;
assign n150 =  ( n32 ) ? ( LB2D_shift_y ) : ( n149 ) ;
assign n151 =  ( n25 ) ? ( n148 ) : ( n150 ) ;
assign n152 =  ( n18 ) ? ( LB2D_shift_y ) : ( n151 ) ;
assign n153 =  ( n9 ) ? ( LB2D_shift_y ) : ( n152 ) ;
assign n154 =  ( n4 ) ? ( LB2D_shift_y ) : ( n153 ) ;
assign n155 =  ( stencil_stream_full ) == ( 1'd1 )  ;
assign n156 =  ( n155 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_0 ) ;
//assign n157 = gb_fun(n156) ;
gb_fun gb_fun_U (
        .stencil (n156),
        .result (n157)
        );

assign n158 =  ( n39 ) ? ( arg_0_TDATA ) : ( arg_0_TDATA ) ;
assign n159 =  ( n32 ) ? ( arg_0_TDATA ) : ( n158 ) ;
assign n160 =  ( n25 ) ? ( arg_0_TDATA ) : ( n159 ) ;
assign n161 =  ( n18 ) ? ( n157 ) : ( n160 ) ;
assign n162 =  ( n9 ) ? ( arg_0_TDATA ) : ( n161 ) ;
assign n163 =  ( n4 ) ? ( arg_0_TDATA ) : ( n162 ) ;
assign n164 =  ( gb_pp_it_8 ) == ( 1'd1 )  ;
assign n165 =  ( n164 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n166 =  ( n39 ) ? ( arg_0_TVALID ) : ( arg_0_TVALID ) ;
assign n167 =  ( n32 ) ? ( arg_0_TVALID ) : ( n166 ) ;
assign n168 =  ( n25 ) ? ( arg_0_TVALID ) : ( n167 ) ;
assign n169 =  ( n18 ) ? ( n165 ) : ( n168 ) ;
assign n170 =  ( n9 ) ? ( arg_0_TVALID ) : ( n169 ) ;
assign n171 =  ( n4 ) ? ( 1'd0 ) : ( n170 ) ;
assign n172 =  ( n39 ) ? ( 1'd1 ) : ( arg_1_TREADY ) ;
assign n173 =  ( n47 ) ? ( 1'd1 ) : ( n172 ) ;
assign n174 =  ( n32 ) ? ( arg_1_TREADY ) : ( n173 ) ;
assign n175 =  ( n25 ) ? ( arg_1_TREADY ) : ( n174 ) ;
assign n176 =  ( n18 ) ? ( arg_1_TREADY ) : ( n175 ) ;
assign n177 =  ( n9 ) ? ( 1'd0 ) : ( n176 ) ;
assign n178 =  ( n4 ) ? ( 1'd0 ) : ( n177 ) ;
assign n179 =  ( gb_p_cnt ) + ( 19'd1 )  ;
assign n180 =  ( n179 ) == ( 19'd307200 )  ;
assign n181 =  ( n180 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n182 =  ( n39 ) ? ( gb_exit_it_1 ) : ( gb_exit_it_1 ) ;
assign n183 =  ( n32 ) ? ( gb_exit_it_1 ) : ( n182 ) ;
assign n184 =  ( n25 ) ? ( gb_exit_it_1 ) : ( n183 ) ;
assign n185 =  ( n18 ) ? ( n181 ) : ( n184 ) ;
assign n186 =  ( n9 ) ? ( gb_exit_it_1 ) : ( n185 ) ;
assign n187 =  ( n4 ) ? ( gb_exit_it_1 ) : ( n186 ) ;
assign n188 =  ( n39 ) ? ( gb_exit_it_2 ) : ( gb_exit_it_2 ) ;
assign n189 =  ( n32 ) ? ( gb_exit_it_2 ) : ( n188 ) ;
assign n190 =  ( n25 ) ? ( gb_exit_it_2 ) : ( n189 ) ;
assign n191 =  ( n18 ) ? ( gb_exit_it_1 ) : ( n190 ) ;
assign n192 =  ( n9 ) ? ( gb_exit_it_2 ) : ( n191 ) ;
assign n193 =  ( n4 ) ? ( gb_exit_it_2 ) : ( n192 ) ;
assign n194 =  ( n39 ) ? ( gb_exit_it_3 ) : ( gb_exit_it_3 ) ;
assign n195 =  ( n32 ) ? ( gb_exit_it_3 ) : ( n194 ) ;
assign n196 =  ( n25 ) ? ( gb_exit_it_3 ) : ( n195 ) ;
assign n197 =  ( n18 ) ? ( gb_exit_it_2 ) : ( n196 ) ;
assign n198 =  ( n9 ) ? ( gb_exit_it_3 ) : ( n197 ) ;
assign n199 =  ( n4 ) ? ( gb_exit_it_3 ) : ( n198 ) ;
assign n200 =  ( n39 ) ? ( gb_exit_it_4 ) : ( gb_exit_it_4 ) ;
assign n201 =  ( n32 ) ? ( gb_exit_it_4 ) : ( n200 ) ;
assign n202 =  ( n25 ) ? ( gb_exit_it_4 ) : ( n201 ) ;
assign n203 =  ( n18 ) ? ( gb_exit_it_3 ) : ( n202 ) ;
assign n204 =  ( n9 ) ? ( gb_exit_it_4 ) : ( n203 ) ;
assign n205 =  ( n4 ) ? ( gb_exit_it_4 ) : ( n204 ) ;
assign n206 =  ( n39 ) ? ( gb_exit_it_5 ) : ( gb_exit_it_5 ) ;
assign n207 =  ( n32 ) ? ( gb_exit_it_5 ) : ( n206 ) ;
assign n208 =  ( n25 ) ? ( gb_exit_it_5 ) : ( n207 ) ;
assign n209 =  ( n18 ) ? ( gb_exit_it_4 ) : ( n208 ) ;
assign n210 =  ( n9 ) ? ( gb_exit_it_5 ) : ( n209 ) ;
assign n211 =  ( n4 ) ? ( gb_exit_it_5 ) : ( n210 ) ;
assign n212 =  ( n39 ) ? ( gb_exit_it_6 ) : ( gb_exit_it_6 ) ;
assign n213 =  ( n32 ) ? ( gb_exit_it_6 ) : ( n212 ) ;
assign n214 =  ( n25 ) ? ( gb_exit_it_6 ) : ( n213 ) ;
assign n215 =  ( n18 ) ? ( gb_exit_it_5 ) : ( n214 ) ;
assign n216 =  ( n9 ) ? ( gb_exit_it_6 ) : ( n215 ) ;
assign n217 =  ( n4 ) ? ( gb_exit_it_6 ) : ( n216 ) ;
assign n218 =  ( n39 ) ? ( gb_exit_it_7 ) : ( gb_exit_it_7 ) ;
assign n219 =  ( n32 ) ? ( gb_exit_it_7 ) : ( n218 ) ;
assign n220 =  ( n25 ) ? ( gb_exit_it_7 ) : ( n219 ) ;
assign n221 =  ( n18 ) ? ( gb_exit_it_6 ) : ( n220 ) ;
assign n222 =  ( n9 ) ? ( gb_exit_it_7 ) : ( n221 ) ;
assign n223 =  ( n4 ) ? ( gb_exit_it_7 ) : ( n222 ) ;
assign n224 =  ( n39 ) ? ( gb_exit_it_8 ) : ( gb_exit_it_8 ) ;
assign n225 =  ( n32 ) ? ( gb_exit_it_8 ) : ( n224 ) ;
assign n226 =  ( n25 ) ? ( gb_exit_it_8 ) : ( n225 ) ;
assign n227 =  ( n18 ) ? ( gb_exit_it_7 ) : ( n226 ) ;
assign n228 =  ( n9 ) ? ( gb_exit_it_8 ) : ( n227 ) ;
assign n229 =  ( n4 ) ? ( gb_exit_it_8 ) : ( n228 ) ;
assign n230 =  ( gb_p_cnt ) < ( 19'd307200 )  ;
assign n231 =  ( n230 ) ? ( n179 ) : ( 19'd307200 ) ;
assign n232 =  ( n39 ) ? ( gb_p_cnt ) : ( gb_p_cnt ) ;
assign n233 =  ( n32 ) ? ( gb_p_cnt ) : ( n232 ) ;
assign n234 =  ( n25 ) ? ( gb_p_cnt ) : ( n233 ) ;
assign n235 =  ( n18 ) ? ( n231 ) : ( n234 ) ;
assign n236 =  ( n9 ) ? ( gb_p_cnt ) : ( n235 ) ;
assign n237 =  ( n4 ) ? ( gb_p_cnt ) : ( n236 ) ;
assign n238 =  ( n39 ) ? ( gb_pp_it_1 ) : ( gb_pp_it_1 ) ;
assign n239 =  ( n32 ) ? ( gb_pp_it_1 ) : ( n238 ) ;
assign n240 =  ( n25 ) ? ( gb_pp_it_1 ) : ( n239 ) ;
assign n241 =  ( n18 ) ? ( 1'd1 ) : ( n240 ) ;
assign n242 =  ( n9 ) ? ( gb_pp_it_1 ) : ( n241 ) ;
assign n243 =  ( n4 ) ? ( gb_pp_it_1 ) : ( n242 ) ;
assign n244 =  ( n39 ) ? ( gb_pp_it_2 ) : ( gb_pp_it_2 ) ;
assign n245 =  ( n32 ) ? ( gb_pp_it_2 ) : ( n244 ) ;
assign n246 =  ( n25 ) ? ( gb_pp_it_2 ) : ( n245 ) ;
assign n247 =  ( n18 ) ? ( gb_pp_it_1 ) : ( n246 ) ;
assign n248 =  ( n9 ) ? ( gb_pp_it_2 ) : ( n247 ) ;
assign n249 =  ( n4 ) ? ( gb_pp_it_2 ) : ( n248 ) ;
assign n250 =  ( n39 ) ? ( gb_pp_it_3 ) : ( gb_pp_it_3 ) ;
assign n251 =  ( n32 ) ? ( gb_pp_it_3 ) : ( n250 ) ;
assign n252 =  ( n25 ) ? ( gb_pp_it_3 ) : ( n251 ) ;
assign n253 =  ( n18 ) ? ( gb_pp_it_2 ) : ( n252 ) ;
assign n254 =  ( n9 ) ? ( gb_pp_it_3 ) : ( n253 ) ;
assign n255 =  ( n4 ) ? ( gb_pp_it_3 ) : ( n254 ) ;
assign n256 =  ( n39 ) ? ( gb_pp_it_4 ) : ( gb_pp_it_4 ) ;
assign n257 =  ( n32 ) ? ( gb_pp_it_4 ) : ( n256 ) ;
assign n258 =  ( n25 ) ? ( gb_pp_it_4 ) : ( n257 ) ;
assign n259 =  ( n18 ) ? ( gb_pp_it_3 ) : ( n258 ) ;
assign n260 =  ( n9 ) ? ( gb_pp_it_4 ) : ( n259 ) ;
assign n261 =  ( n4 ) ? ( gb_pp_it_4 ) : ( n260 ) ;
assign n262 =  ( n39 ) ? ( gb_pp_it_5 ) : ( gb_pp_it_5 ) ;
assign n263 =  ( n32 ) ? ( gb_pp_it_5 ) : ( n262 ) ;
assign n264 =  ( n25 ) ? ( gb_pp_it_5 ) : ( n263 ) ;
assign n265 =  ( n18 ) ? ( gb_pp_it_4 ) : ( n264 ) ;
assign n266 =  ( n9 ) ? ( gb_pp_it_5 ) : ( n265 ) ;
assign n267 =  ( n4 ) ? ( gb_pp_it_5 ) : ( n266 ) ;
assign n268 =  ( n39 ) ? ( gb_pp_it_6 ) : ( gb_pp_it_6 ) ;
assign n269 =  ( n32 ) ? ( gb_pp_it_6 ) : ( n268 ) ;
assign n270 =  ( n25 ) ? ( gb_pp_it_6 ) : ( n269 ) ;
assign n271 =  ( n18 ) ? ( gb_pp_it_5 ) : ( n270 ) ;
assign n272 =  ( n9 ) ? ( gb_pp_it_6 ) : ( n271 ) ;
assign n273 =  ( n4 ) ? ( gb_pp_it_6 ) : ( n272 ) ;
assign n274 =  ( n39 ) ? ( gb_pp_it_7 ) : ( gb_pp_it_7 ) ;
assign n275 =  ( n32 ) ? ( gb_pp_it_7 ) : ( n274 ) ;
assign n276 =  ( n25 ) ? ( gb_pp_it_7 ) : ( n275 ) ;
assign n277 =  ( n18 ) ? ( gb_pp_it_6 ) : ( n276 ) ;
assign n278 =  ( n9 ) ? ( gb_pp_it_7 ) : ( n277 ) ;
assign n279 =  ( n4 ) ? ( gb_pp_it_7 ) : ( n278 ) ;
assign n280 =  ( n39 ) ? ( gb_pp_it_8 ) : ( gb_pp_it_8 ) ;
assign n281 =  ( n32 ) ? ( gb_pp_it_8 ) : ( n280 ) ;
assign n282 =  ( n25 ) ? ( gb_pp_it_8 ) : ( n281 ) ;
assign n283 =  ( n18 ) ? ( gb_pp_it_7 ) : ( n282 ) ;
assign n284 =  ( n9 ) ? ( gb_pp_it_8 ) : ( n283 ) ;
assign n285 =  ( n4 ) ? ( gb_pp_it_8 ) : ( n284 ) ;
assign n286 =  ( n39 ) ? ( gb_pp_it_9 ) : ( gb_pp_it_9 ) ;
assign n287 =  ( n32 ) ? ( gb_pp_it_9 ) : ( n286 ) ;
assign n288 =  ( n25 ) ? ( gb_pp_it_9 ) : ( n287 ) ;
assign n289 =  ( n18 ) ? ( gb_pp_it_8 ) : ( n288 ) ;
assign n290 =  ( n9 ) ? ( gb_pp_it_9 ) : ( n289 ) ;
assign n291 =  ( n4 ) ? ( gb_pp_it_9 ) : ( n290 ) ;
assign n292 =  ( n39 ) ? ( LB1D_buff ) : ( in_stream_buff_0 ) ;
assign n293 =  ( n32 ) ? ( in_stream_buff_0 ) : ( n292 ) ;
assign n294 =  ( n25 ) ? ( in_stream_buff_0 ) : ( n293 ) ;
assign n295 =  ( n18 ) ? ( in_stream_buff_0 ) : ( n294 ) ;
assign n296 =  ( n9 ) ? ( in_stream_buff_0 ) : ( n295 ) ;
assign n297 =  ( n4 ) ? ( in_stream_buff_0 ) : ( n296 ) ;
assign n298 =  ( n39 ) ? ( in_stream_buff_0 ) : ( in_stream_buff_1 ) ;
assign n299 =  ( n32 ) ? ( in_stream_buff_1 ) : ( n298 ) ;
assign n300 =  ( n25 ) ? ( in_stream_buff_1 ) : ( n299 ) ;
assign n301 =  ( n18 ) ? ( in_stream_buff_1 ) : ( n300 ) ;
assign n302 =  ( n9 ) ? ( in_stream_buff_1 ) : ( n301 ) ;
assign n303 =  ( n4 ) ? ( in_stream_buff_1 ) : ( n302 ) ;
assign n304 =  ( in_stream_full ) == ( 1'd1 )  ;
assign n305 =  ( n304 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n306 =  ( n39 ) ? ( 1'd0 ) : ( in_stream_empty ) ;
assign n307 =  ( n32 ) ? ( n305 ) : ( n306 ) ;
assign n308 =  ( n25 ) ? ( in_stream_empty ) : ( n307 ) ;
assign n309 =  ( n18 ) ? ( in_stream_empty ) : ( n308 ) ;
assign n310 =  ( n9 ) ? ( in_stream_empty ) : ( n309 ) ;
assign n311 =  ( n4 ) ? ( in_stream_empty ) : ( n310 ) ;
assign n312 =  ( in_stream_empty ) == ( 1'd1 )  ;
assign n313 =  ( n312 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n314 =  ( n39 ) ? ( n313 ) : ( in_stream_full ) ;
assign n315 =  ( n32 ) ? ( 1'd0 ) : ( n314 ) ;
assign n316 =  ( n25 ) ? ( in_stream_full ) : ( n315 ) ;
assign n317 =  ( n18 ) ? ( in_stream_full ) : ( n316 ) ;
assign n318 =  ( n9 ) ? ( in_stream_full ) : ( n317 ) ;
assign n319 =  ( n4 ) ? ( in_stream_full ) : ( n318 ) ;
assign n320 =  ( n304 ) ? ( in_stream_buff_1 ) : ( in_stream_buff_0 ) ;
assign n321 =  ( LB2D_proc_w ) == ( 64'd0 )  ;
assign n322 =  (  LB2D_proc_7 [ LB2D_proc_x ] )  ;
assign n323 =  ( LB2D_proc_w ) == ( 64'd1 )  ;
assign n324 =  (  LB2D_proc_0 [ LB2D_proc_x ] )  ;
assign n325 =  ( LB2D_proc_w ) == ( 64'd2 )  ;
assign n326 =  (  LB2D_proc_1 [ LB2D_proc_x ] )  ;
assign n327 =  ( LB2D_proc_w ) == ( 64'd3 )  ;
assign n328 =  (  LB2D_proc_2 [ LB2D_proc_x ] )  ;
assign n329 =  ( LB2D_proc_w ) == ( 64'd4 )  ;
assign n330 =  (  LB2D_proc_3 [ LB2D_proc_x ] )  ;
assign n331 =  ( LB2D_proc_w ) == ( 64'd5 )  ;
assign n332 =  (  LB2D_proc_4 [ LB2D_proc_x ] )  ;
assign n333 =  ( LB2D_proc_w ) == ( 64'd6 )  ;
assign n334 =  (  LB2D_proc_5 [ LB2D_proc_x ] )  ;
assign n335 =  (  LB2D_proc_6 [ LB2D_proc_x ] )  ;
assign n336 =  ( n333 ) ? ( n334 ) : ( n335 ) ;
assign n337 =  ( n331 ) ? ( n332 ) : ( n336 ) ;
assign n338 =  ( n329 ) ? ( n330 ) : ( n337 ) ;
assign n339 =  ( n327 ) ? ( n328 ) : ( n338 ) ;
assign n340 =  ( n325 ) ? ( n326 ) : ( n339 ) ;
assign n341 =  ( n323 ) ? ( n324 ) : ( n340 ) ;
assign n342 =  ( n321 ) ? ( n322 ) : ( n341 ) ;
assign n343 =  ( n333 ) ? ( n332 ) : ( n334 ) ;
assign n344 =  ( n331 ) ? ( n330 ) : ( n343 ) ;
assign n345 =  ( n329 ) ? ( n328 ) : ( n344 ) ;
assign n346 =  ( n327 ) ? ( n326 ) : ( n345 ) ;
assign n347 =  ( n325 ) ? ( n324 ) : ( n346 ) ;
assign n348 =  ( n323 ) ? ( n322 ) : ( n347 ) ;
assign n349 =  ( n321 ) ? ( n335 ) : ( n348 ) ;
assign n350 =  ( n333 ) ? ( n330 ) : ( n332 ) ;
assign n351 =  ( n331 ) ? ( n328 ) : ( n350 ) ;
assign n352 =  ( n329 ) ? ( n326 ) : ( n351 ) ;
assign n353 =  ( n327 ) ? ( n324 ) : ( n352 ) ;
assign n354 =  ( n325 ) ? ( n322 ) : ( n353 ) ;
assign n355 =  ( n323 ) ? ( n335 ) : ( n354 ) ;
assign n356 =  ( n321 ) ? ( n334 ) : ( n355 ) ;
assign n357 =  ( n333 ) ? ( n328 ) : ( n330 ) ;
assign n358 =  ( n331 ) ? ( n326 ) : ( n357 ) ;
assign n359 =  ( n329 ) ? ( n324 ) : ( n358 ) ;
assign n360 =  ( n327 ) ? ( n322 ) : ( n359 ) ;
assign n361 =  ( n325 ) ? ( n335 ) : ( n360 ) ;
assign n362 =  ( n323 ) ? ( n334 ) : ( n361 ) ;
assign n363 =  ( n321 ) ? ( n332 ) : ( n362 ) ;
assign n364 =  ( n333 ) ? ( n326 ) : ( n328 ) ;
assign n365 =  ( n331 ) ? ( n324 ) : ( n364 ) ;
assign n366 =  ( n329 ) ? ( n322 ) : ( n365 ) ;
assign n367 =  ( n327 ) ? ( n335 ) : ( n366 ) ;
assign n368 =  ( n325 ) ? ( n334 ) : ( n367 ) ;
assign n369 =  ( n323 ) ? ( n332 ) : ( n368 ) ;
assign n370 =  ( n321 ) ? ( n330 ) : ( n369 ) ;
assign n371 =  ( n333 ) ? ( n324 ) : ( n326 ) ;
assign n372 =  ( n331 ) ? ( n322 ) : ( n371 ) ;
assign n373 =  ( n329 ) ? ( n335 ) : ( n372 ) ;
assign n374 =  ( n327 ) ? ( n334 ) : ( n373 ) ;
assign n375 =  ( n325 ) ? ( n332 ) : ( n374 ) ;
assign n376 =  ( n323 ) ? ( n330 ) : ( n375 ) ;
assign n377 =  ( n321 ) ? ( n328 ) : ( n376 ) ;
assign n378 =  ( n333 ) ? ( n322 ) : ( n324 ) ;
assign n379 =  ( n331 ) ? ( n335 ) : ( n378 ) ;
assign n380 =  ( n329 ) ? ( n334 ) : ( n379 ) ;
assign n381 =  ( n327 ) ? ( n332 ) : ( n380 ) ;
assign n382 =  ( n325 ) ? ( n330 ) : ( n381 ) ;
assign n383 =  ( n323 ) ? ( n328 ) : ( n382 ) ;
assign n384 =  ( n321 ) ? ( n326 ) : ( n383 ) ;
assign n385 =  ( n333 ) ? ( n335 ) : ( n322 ) ;
assign n386 =  ( n331 ) ? ( n334 ) : ( n385 ) ;
assign n387 =  ( n329 ) ? ( n332 ) : ( n386 ) ;
assign n388 =  ( n327 ) ? ( n330 ) : ( n387 ) ;
assign n389 =  ( n325 ) ? ( n328 ) : ( n388 ) ;
assign n390 =  ( n323 ) ? ( n326 ) : ( n389 ) ;
assign n391 =  ( n321 ) ? ( n324 ) : ( n390 ) ;
assign n392 =  { ( n384 ) , ( n391 ) }  ;
assign n393 =  { ( n377 ) , ( n392 ) }  ;
assign n394 =  { ( n370 ) , ( n393 ) }  ;
assign n395 =  { ( n363 ) , ( n394 ) }  ;
assign n396 =  { ( n356 ) , ( n395 ) }  ;
assign n397 =  { ( n349 ) , ( n396 ) }  ;
assign n398 =  { ( n342 ) , ( n397 ) }  ;
assign n399 =  { ( n320 ) , ( n398 ) }  ;
assign n400 =  ( n30 ) ? ( slice_stream_buff_0 ) : ( n399 ) ;
assign n401 =  ( n39 ) ? ( slice_stream_buff_0 ) : ( slice_stream_buff_0 ) ;
assign n402 =  ( n32 ) ? ( n400 ) : ( n401 ) ;
assign n403 =  ( n25 ) ? ( slice_stream_buff_0 ) : ( n402 ) ;
assign n404 =  ( n18 ) ? ( slice_stream_buff_0 ) : ( n403 ) ;
assign n405 =  ( n9 ) ? ( slice_stream_buff_0 ) : ( n404 ) ;
assign n406 =  ( n4 ) ? ( slice_stream_buff_0 ) : ( n405 ) ;
assign n407 =  ( n30 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n408 =  ( n39 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_1 ) ;
assign n409 =  ( n32 ) ? ( n407 ) : ( n408 ) ;
assign n410 =  ( n25 ) ? ( slice_stream_buff_1 ) : ( n409 ) ;
assign n411 =  ( n18 ) ? ( slice_stream_buff_1 ) : ( n410 ) ;
assign n412 =  ( n9 ) ? ( slice_stream_buff_1 ) : ( n411 ) ;
assign n413 =  ( n4 ) ? ( slice_stream_buff_1 ) : ( n412 ) ;
assign n414 =  ( n87 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n415 =  ( n30 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n416 =  ( n39 ) ? ( slice_stream_empty ) : ( slice_stream_empty ) ;
assign n417 =  ( n32 ) ? ( n415 ) : ( n416 ) ;
assign n418 =  ( n25 ) ? ( n414 ) : ( n417 ) ;
assign n419 =  ( n18 ) ? ( slice_stream_empty ) : ( n418 ) ;
assign n420 =  ( n9 ) ? ( slice_stream_empty ) : ( n419 ) ;
assign n421 =  ( n4 ) ? ( slice_stream_empty ) : ( n420 ) ;
assign n422 =  ( slice_stream_empty ) == ( 1'd1 )  ;
assign n423 =  ( n422 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n424 =  ( n30 ) ? ( 1'd0 ) : ( n423 ) ;
assign n425 =  ( n39 ) ? ( slice_stream_full ) : ( slice_stream_full ) ;
assign n426 =  ( n32 ) ? ( n424 ) : ( n425 ) ;
assign n427 =  ( n25 ) ? ( 1'd0 ) : ( n426 ) ;
assign n428 =  ( n18 ) ? ( slice_stream_full ) : ( n427 ) ;
assign n429 =  ( n9 ) ? ( slice_stream_full ) : ( n428 ) ;
assign n430 =  ( n4 ) ? ( slice_stream_full ) : ( n429 ) ;
assign n431 =  ( LB2D_shift_x ) >= ( 9'd8 )  ;
assign n432 = n88[71:64] ;
assign n433 = LB2D_shift_0[71:64] ;
assign n434 = LB2D_shift_1[71:64] ;
assign n435 = LB2D_shift_2[71:64] ;
assign n436 = LB2D_shift_3[71:64] ;
assign n437 = LB2D_shift_4[71:64] ;
assign n438 = LB2D_shift_5[71:64] ;
assign n439 = LB2D_shift_6[71:64] ;
assign n440 = LB2D_shift_7[71:64] ;
assign n441 =  { ( n439 ) , ( n440 ) }  ;
assign n442 =  { ( n438 ) , ( n441 ) }  ;
assign n443 =  { ( n437 ) , ( n442 ) }  ;
assign n444 =  { ( n436 ) , ( n443 ) }  ;
assign n445 =  { ( n435 ) , ( n444 ) }  ;
assign n446 =  { ( n434 ) , ( n445 ) }  ;
assign n447 =  { ( n433 ) , ( n446 ) }  ;
assign n448 =  { ( n432 ) , ( n447 ) }  ;
assign n449 = n88[63:56] ;
assign n450 = LB2D_shift_0[63:56] ;
assign n451 = LB2D_shift_1[63:56] ;
assign n452 = LB2D_shift_2[63:56] ;
assign n453 = LB2D_shift_3[63:56] ;
assign n454 = LB2D_shift_4[63:56] ;
assign n455 = LB2D_shift_5[63:56] ;
assign n456 = LB2D_shift_6[63:56] ;
assign n457 = LB2D_shift_7[63:56] ;
assign n458 =  { ( n456 ) , ( n457 ) }  ;
assign n459 =  { ( n455 ) , ( n458 ) }  ;
assign n460 =  { ( n454 ) , ( n459 ) }  ;
assign n461 =  { ( n453 ) , ( n460 ) }  ;
assign n462 =  { ( n452 ) , ( n461 ) }  ;
assign n463 =  { ( n451 ) , ( n462 ) }  ;
assign n464 =  { ( n450 ) , ( n463 ) }  ;
assign n465 =  { ( n449 ) , ( n464 ) }  ;
assign n466 = n88[55:48] ;
assign n467 = LB2D_shift_0[55:48] ;
assign n468 = LB2D_shift_1[55:48] ;
assign n469 = LB2D_shift_2[55:48] ;
assign n470 = LB2D_shift_3[55:48] ;
assign n471 = LB2D_shift_4[55:48] ;
assign n472 = LB2D_shift_5[55:48] ;
assign n473 = LB2D_shift_6[55:48] ;
assign n474 = LB2D_shift_7[55:48] ;
assign n475 =  { ( n473 ) , ( n474 ) }  ;
assign n476 =  { ( n472 ) , ( n475 ) }  ;
assign n477 =  { ( n471 ) , ( n476 ) }  ;
assign n478 =  { ( n470 ) , ( n477 ) }  ;
assign n479 =  { ( n469 ) , ( n478 ) }  ;
assign n480 =  { ( n468 ) , ( n479 ) }  ;
assign n481 =  { ( n467 ) , ( n480 ) }  ;
assign n482 =  { ( n466 ) , ( n481 ) }  ;
assign n483 = n88[47:40] ;
assign n484 = LB2D_shift_0[47:40] ;
assign n485 = LB2D_shift_1[47:40] ;
assign n486 = LB2D_shift_2[47:40] ;
assign n487 = LB2D_shift_3[47:40] ;
assign n488 = LB2D_shift_4[47:40] ;
assign n489 = LB2D_shift_5[47:40] ;
assign n490 = LB2D_shift_6[47:40] ;
assign n491 = LB2D_shift_7[47:40] ;
assign n492 =  { ( n490 ) , ( n491 ) }  ;
assign n493 =  { ( n489 ) , ( n492 ) }  ;
assign n494 =  { ( n488 ) , ( n493 ) }  ;
assign n495 =  { ( n487 ) , ( n494 ) }  ;
assign n496 =  { ( n486 ) , ( n495 ) }  ;
assign n497 =  { ( n485 ) , ( n496 ) }  ;
assign n498 =  { ( n484 ) , ( n497 ) }  ;
assign n499 =  { ( n483 ) , ( n498 ) }  ;
assign n500 = n88[39:32] ;
assign n501 = LB2D_shift_0[39:32] ;
assign n502 = LB2D_shift_1[39:32] ;
assign n503 = LB2D_shift_2[39:32] ;
assign n504 = LB2D_shift_3[39:32] ;
assign n505 = LB2D_shift_4[39:32] ;
assign n506 = LB2D_shift_5[39:32] ;
assign n507 = LB2D_shift_6[39:32] ;
assign n508 = LB2D_shift_7[39:32] ;
assign n509 =  { ( n507 ) , ( n508 ) }  ;
assign n510 =  { ( n506 ) , ( n509 ) }  ;
assign n511 =  { ( n505 ) , ( n510 ) }  ;
assign n512 =  { ( n504 ) , ( n511 ) }  ;
assign n513 =  { ( n503 ) , ( n512 ) }  ;
assign n514 =  { ( n502 ) , ( n513 ) }  ;
assign n515 =  { ( n501 ) , ( n514 ) }  ;
assign n516 =  { ( n500 ) , ( n515 ) }  ;
assign n517 = n88[31:24] ;
assign n518 = LB2D_shift_0[31:24] ;
assign n519 = LB2D_shift_1[31:24] ;
assign n520 = LB2D_shift_2[31:24] ;
assign n521 = LB2D_shift_3[31:24] ;
assign n522 = LB2D_shift_4[31:24] ;
assign n523 = LB2D_shift_5[31:24] ;
assign n524 = LB2D_shift_6[31:24] ;
assign n525 = LB2D_shift_7[31:24] ;
assign n526 =  { ( n524 ) , ( n525 ) }  ;
assign n527 =  { ( n523 ) , ( n526 ) }  ;
assign n528 =  { ( n522 ) , ( n527 ) }  ;
assign n529 =  { ( n521 ) , ( n528 ) }  ;
assign n530 =  { ( n520 ) , ( n529 ) }  ;
assign n531 =  { ( n519 ) , ( n530 ) }  ;
assign n532 =  { ( n518 ) , ( n531 ) }  ;
assign n533 =  { ( n517 ) , ( n532 ) }  ;
assign n534 = n88[23:16] ;
assign n535 = LB2D_shift_0[23:16] ;
assign n536 = LB2D_shift_1[23:16] ;
assign n537 = LB2D_shift_2[23:16] ;
assign n538 = LB2D_shift_3[23:16] ;
assign n539 = LB2D_shift_4[23:16] ;
assign n540 = LB2D_shift_5[23:16] ;
assign n541 = LB2D_shift_6[23:16] ;
assign n542 = LB2D_shift_7[23:16] ;
assign n543 =  { ( n541 ) , ( n542 ) }  ;
assign n544 =  { ( n540 ) , ( n543 ) }  ;
assign n545 =  { ( n539 ) , ( n544 ) }  ;
assign n546 =  { ( n538 ) , ( n545 ) }  ;
assign n547 =  { ( n537 ) , ( n546 ) }  ;
assign n548 =  { ( n536 ) , ( n547 ) }  ;
assign n549 =  { ( n535 ) , ( n548 ) }  ;
assign n550 =  { ( n534 ) , ( n549 ) }  ;
assign n551 = n88[15:8] ;
assign n552 = LB2D_shift_0[15:8] ;
assign n553 = LB2D_shift_1[15:8] ;
assign n554 = LB2D_shift_2[15:8] ;
assign n555 = LB2D_shift_3[15:8] ;
assign n556 = LB2D_shift_4[15:8] ;
assign n557 = LB2D_shift_5[15:8] ;
assign n558 = LB2D_shift_6[15:8] ;
assign n559 = LB2D_shift_7[15:8] ;
assign n560 =  { ( n558 ) , ( n559 ) }  ;
assign n561 =  { ( n557 ) , ( n560 ) }  ;
assign n562 =  { ( n556 ) , ( n561 ) }  ;
assign n563 =  { ( n555 ) , ( n562 ) }  ;
assign n564 =  { ( n554 ) , ( n563 ) }  ;
assign n565 =  { ( n553 ) , ( n564 ) }  ;
assign n566 =  { ( n552 ) , ( n565 ) }  ;
assign n567 =  { ( n551 ) , ( n566 ) }  ;
assign n568 = n88[7:0] ;
assign n569 = LB2D_shift_0[7:0] ;
assign n570 = LB2D_shift_1[7:0] ;
assign n571 = LB2D_shift_2[7:0] ;
assign n572 = LB2D_shift_3[7:0] ;
assign n573 = LB2D_shift_4[7:0] ;
assign n574 = LB2D_shift_5[7:0] ;
assign n575 = LB2D_shift_6[7:0] ;
assign n576 = LB2D_shift_7[7:0] ;
assign n577 =  { ( n575 ) , ( n576 ) }  ;
assign n578 =  { ( n574 ) , ( n577 ) }  ;
assign n579 =  { ( n573 ) , ( n578 ) }  ;
assign n580 =  { ( n572 ) , ( n579 ) }  ;
assign n581 =  { ( n571 ) , ( n580 ) }  ;
assign n582 =  { ( n570 ) , ( n581 ) }  ;
assign n583 =  { ( n569 ) , ( n582 ) }  ;
assign n584 =  { ( n568 ) , ( n583 ) }  ;
assign n585 =  { ( n567 ) , ( n584 ) }  ;
assign n586 =  { ( n550 ) , ( n585 ) }  ;
assign n587 =  { ( n533 ) , ( n586 ) }  ;
assign n588 =  { ( n516 ) , ( n587 ) }  ;
assign n589 =  { ( n499 ) , ( n588 ) }  ;
assign n590 =  { ( n482 ) , ( n589 ) }  ;
assign n591 =  { ( n465 ) , ( n590 ) }  ;
assign n592 =  { ( n448 ) , ( n591 ) }  ;
assign n593 =  ( n431 ) ? ( n592 ) : ( stencil_stream_buff_0 ) ;
assign n594 =  ( n39 ) ? ( stencil_stream_buff_0 ) : ( stencil_stream_buff_0 ) ;
assign n595 =  ( n32 ) ? ( stencil_stream_buff_0 ) : ( n594 ) ;
assign n596 =  ( n25 ) ? ( n593 ) : ( n595 ) ;
assign n597 =  ( n18 ) ? ( stencil_stream_buff_0 ) : ( n596 ) ;
assign n598 =  ( n9 ) ? ( stencil_stream_buff_0 ) : ( n597 ) ;
assign n599 =  ( n4 ) ? ( stencil_stream_buff_0 ) : ( n598 ) ;
assign n600 =  ( n39 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_1 ) ;
assign n601 =  ( n32 ) ? ( stencil_stream_buff_1 ) : ( n600 ) ;
assign n602 =  ( n25 ) ? ( stencil_stream_buff_0 ) : ( n601 ) ;
assign n603 =  ( n18 ) ? ( stencil_stream_buff_1 ) : ( n602 ) ;
assign n604 =  ( n9 ) ? ( stencil_stream_buff_1 ) : ( n603 ) ;
assign n605 =  ( n4 ) ? ( stencil_stream_buff_1 ) : ( n604 ) ;
assign n606 =  ( n155 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n607 =  ( n23 ) ? ( stencil_stream_empty ) : ( 1'd0 ) ;
assign n608 =  ( n39 ) ? ( stencil_stream_empty ) : ( stencil_stream_empty ) ;
assign n609 =  ( n32 ) ? ( stencil_stream_empty ) : ( n608 ) ;
assign n610 =  ( n25 ) ? ( n607 ) : ( n609 ) ;
assign n611 =  ( n18 ) ? ( n606 ) : ( n610 ) ;
assign n612 =  ( n9 ) ? ( stencil_stream_empty ) : ( n611 ) ;
assign n613 =  ( n4 ) ? ( stencil_stream_empty ) : ( n612 ) ;
assign n614 =  ( n14 ) ? ( 1'd0 ) : ( 1'd0 ) ;
assign n615 =  ( stencil_stream_empty ) == ( 1'd1 )  ;
assign n616 =  ( n615 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n617 =  ( n23 ) ? ( stencil_stream_full ) : ( n616 ) ;
assign n618 =  ( n39 ) ? ( stencil_stream_full ) : ( stencil_stream_full ) ;
assign n619 =  ( n32 ) ? ( stencil_stream_full ) : ( n618 ) ;
assign n620 =  ( n25 ) ? ( n617 ) : ( n619 ) ;
assign n621 =  ( n18 ) ? ( n614 ) : ( n620 ) ;
assign n622 =  ( n9 ) ? ( stencil_stream_full ) : ( n621 ) ;
assign n623 =  ( n4 ) ? ( stencil_stream_full ) : ( n622 ) ;
assign n624 = ~ ( n4 ) ;
assign n625 = ~ ( n9 ) ;
assign n626 =  ( n624 ) & ( n625 )  ;
assign n627 = ~ ( n18 ) ;
assign n628 =  ( n626 ) & ( n627 )  ;
assign n629 = ~ ( n25 ) ;
assign n630 =  ( n628 ) & ( n629 )  ;
assign n631 = ~ ( n32 ) ;
assign n632 =  ( n630 ) & ( n631 )  ;
assign n633 = ~ ( n39 ) ;
assign n634 =  ( n632 ) & ( n633 )  ;
assign n635 =  ( n632 ) & ( n39 )  ;
assign n636 =  ( n630 ) & ( n32 )  ;
assign n637 = ~ ( n321 ) ;
assign n638 =  ( n636 ) & ( n637 )  ;
assign n639 =  ( n636 ) & ( n321 )  ;
assign n640 =  ( n628 ) & ( n25 )  ;
assign n641 =  ( n626 ) & ( n18 )  ;
assign n642 =  ( n624 ) & ( n9 )  ;
assign LB2D_proc_0_addr0 = n639 ? (LB2D_proc_x) : (0);
assign LB2D_proc_0_data0 = n639 ? (n320) : (LB2D_proc_0[0]);
assign n643 = ~ ( n323 ) ;
assign n644 =  ( n636 ) & ( n643 )  ;
assign n645 =  ( n636 ) & ( n323 )  ;
assign LB2D_proc_1_addr0 = n645 ? (LB2D_proc_x) : (0);
assign LB2D_proc_1_data0 = n645 ? (n320) : (LB2D_proc_1[0]);
assign n646 = ~ ( n325 ) ;
assign n647 =  ( n636 ) & ( n646 )  ;
assign n648 =  ( n636 ) & ( n325 )  ;
assign LB2D_proc_2_addr0 = n648 ? (LB2D_proc_x) : (0);
assign LB2D_proc_2_data0 = n648 ? (n320) : (LB2D_proc_2[0]);
assign n649 = ~ ( n327 ) ;
assign n650 =  ( n636 ) & ( n649 )  ;
assign n651 =  ( n636 ) & ( n327 )  ;
assign LB2D_proc_3_addr0 = n651 ? (LB2D_proc_x) : (0);
assign LB2D_proc_3_data0 = n651 ? (n320) : (LB2D_proc_3[0]);
assign n652 = ~ ( n329 ) ;
assign n653 =  ( n636 ) & ( n652 )  ;
assign n654 =  ( n636 ) & ( n329 )  ;
assign LB2D_proc_4_addr0 = n654 ? (LB2D_proc_x) : (0);
assign LB2D_proc_4_data0 = n654 ? (n320) : (LB2D_proc_4[0]);
assign n655 = ~ ( n331 ) ;
assign n656 =  ( n636 ) & ( n655 )  ;
assign n657 =  ( n636 ) & ( n331 )  ;
assign LB2D_proc_5_addr0 = n657 ? (LB2D_proc_x) : (0);
assign LB2D_proc_5_data0 = n657 ? (n320) : (LB2D_proc_5[0]);
assign n658 = ~ ( n333 ) ;
assign n659 =  ( n636 ) & ( n658 )  ;
assign n660 =  ( n636 ) & ( n333 )  ;
assign LB2D_proc_6_addr0 = n660 ? (LB2D_proc_x) : (0);
assign LB2D_proc_6_data0 = n660 ? (n320) : (LB2D_proc_6[0]);
assign n661 =  ( LB2D_proc_w ) == ( 64'd7 )  ;
assign n662 = ~ ( n661 ) ;
assign n663 =  ( n636 ) & ( n662 )  ;
assign n664 =  ( n636 ) & ( n661 )  ;
assign LB2D_proc_7_addr0 = n664 ? (LB2D_proc_x) : (0);
assign LB2D_proc_7_data0 = n664 ? (n320) : (LB2D_proc_7[0]);
/*
function [7:0] gb_fun ;
input [647:0] arg0;
    begin
//TODO: Add the specific function HERE.    end
endfunction
*/

always @(posedge clk) begin
   if(rst) begin
       LB1D_buff <= LB1D_buff;
       LB1D_it_1 <= LB1D_it_1;
       LB1D_p_cnt <= LB1D_p_cnt;
       LB2D_proc_w <= LB2D_proc_w;
       LB2D_proc_x <= LB2D_proc_x;
       LB2D_proc_y <= LB2D_proc_y;
       LB2D_shift_0 <= LB2D_shift_0;
       LB2D_shift_1 <= LB2D_shift_1;
       LB2D_shift_2 <= LB2D_shift_2;
       LB2D_shift_3 <= LB2D_shift_3;
       LB2D_shift_4 <= LB2D_shift_4;
       LB2D_shift_5 <= LB2D_shift_5;
       LB2D_shift_6 <= LB2D_shift_6;
       LB2D_shift_7 <= LB2D_shift_7;
       LB2D_shift_x <= LB2D_shift_x;
       LB2D_shift_y <= LB2D_shift_y;
       arg_0_TDATA <= arg_0_TDATA;
       arg_0_TVALID <= arg_0_TVALID;
       arg_1_TREADY <= arg_1_TREADY;
       gb_exit_it_1 <= gb_exit_it_1;
       gb_exit_it_2 <= gb_exit_it_2;
       gb_exit_it_3 <= gb_exit_it_3;
       gb_exit_it_4 <= gb_exit_it_4;
       gb_exit_it_5 <= gb_exit_it_5;
       gb_exit_it_6 <= gb_exit_it_6;
       gb_exit_it_7 <= gb_exit_it_7;
       gb_exit_it_8 <= gb_exit_it_8;
       gb_p_cnt <= gb_p_cnt;
       gb_pp_it_1 <= gb_pp_it_1;
       gb_pp_it_2 <= gb_pp_it_2;
       gb_pp_it_3 <= gb_pp_it_3;
       gb_pp_it_4 <= gb_pp_it_4;
       gb_pp_it_5 <= gb_pp_it_5;
       gb_pp_it_6 <= gb_pp_it_6;
       gb_pp_it_7 <= gb_pp_it_7;
       gb_pp_it_8 <= gb_pp_it_8;
       gb_pp_it_9 <= gb_pp_it_9;
       in_stream_buff_0 <= in_stream_buff_0;
       in_stream_buff_1 <= in_stream_buff_1;
       in_stream_empty <= in_stream_empty;
       in_stream_full <= in_stream_full;
       slice_stream_buff_0 <= slice_stream_buff_0;
       slice_stream_buff_1 <= slice_stream_buff_1;
       slice_stream_empty <= slice_stream_empty;
       slice_stream_full <= slice_stream_full;
       stencil_stream_buff_0 <= stencil_stream_buff_0;
       stencil_stream_buff_1 <= stencil_stream_buff_1;
       stencil_stream_empty <= stencil_stream_empty;
       stencil_stream_full <= stencil_stream_full;
   end
   else if(step) begin
       LB1D_buff <= n45;
       LB1D_it_1 <= n48;
       LB1D_p_cnt <= n56;
       LB2D_proc_w <= n67;
       LB2D_proc_x <= n78;
       LB2D_proc_y <= n86;
       LB2D_shift_0 <= n94;
       LB2D_shift_1 <= n100;
       LB2D_shift_2 <= n106;
       LB2D_shift_3 <= n112;
       LB2D_shift_4 <= n118;
       LB2D_shift_5 <= n124;
       LB2D_shift_6 <= n130;
       LB2D_shift_7 <= n136;
       LB2D_shift_x <= n143;
       LB2D_shift_y <= n154;
       arg_0_TDATA <= n163;
       arg_0_TVALID <= n171;
       arg_1_TREADY <= n178;
       gb_exit_it_1 <= n187;
       gb_exit_it_2 <= n193;
       gb_exit_it_3 <= n199;
       gb_exit_it_4 <= n205;
       gb_exit_it_5 <= n211;
       gb_exit_it_6 <= n217;
       gb_exit_it_7 <= n223;
       gb_exit_it_8 <= n229;
       gb_p_cnt <= n237;
       gb_pp_it_1 <= n243;
       gb_pp_it_2 <= n249;
       gb_pp_it_3 <= n255;
       gb_pp_it_4 <= n261;
       gb_pp_it_5 <= n267;
       gb_pp_it_6 <= n273;
       gb_pp_it_7 <= n279;
       gb_pp_it_8 <= n285;
       gb_pp_it_9 <= n291;
       in_stream_buff_0 <= n297;
       in_stream_buff_1 <= n303;
       in_stream_empty <= n311;
       in_stream_full <= n319;
       slice_stream_buff_0 <= n406;
       slice_stream_buff_1 <= n413;
       slice_stream_empty <= n421;
       slice_stream_full <= n430;
       stencil_stream_buff_0 <= n599;
       stencil_stream_buff_1 <= n605;
       stencil_stream_empty <= n613;
       stencil_stream_full <= n623;
       LB2D_proc_0 [ LB2D_proc_0_addr0 ] <= LB2D_proc_0_data0;
       LB2D_proc_1 [ LB2D_proc_1_addr0 ] <= LB2D_proc_1_data0;
       LB2D_proc_2 [ LB2D_proc_2_addr0 ] <= LB2D_proc_2_data0;
       LB2D_proc_3 [ LB2D_proc_3_addr0 ] <= LB2D_proc_3_data0;
       LB2D_proc_4 [ LB2D_proc_4_addr0 ] <= LB2D_proc_4_data0;
       LB2D_proc_5 [ LB2D_proc_5_addr0 ] <= LB2D_proc_5_data0;
       LB2D_proc_6 [ LB2D_proc_6_addr0 ] <= LB2D_proc_6_data0;
       LB2D_proc_7 [ LB2D_proc_7_addr0 ] <= LB2D_proc_7_data0;
   end
end
endmodule
