module GB(
arg_0_TREADY,
arg_1_TDATA,
arg_1_TVALID,
LB1D_buff,
LB2D_proc_w,
LB2D_proc_x,
LB2D_proc_y,
LB2D_shift_0,
LB2D_shift_1,
LB2D_shift_2,
LB2D_shift_3,
LB2D_shift_4,
LB2D_shift_5,
LB2D_shift_6,
LB2D_shift_7,
LB2D_shift_x,
LB2D_shift_y,
arg_0_TDATA,
arg_0_TVALID,
arg_1_TREADY,
in_stream_buff_0,
in_stream_buff_1,
in_stream_empty,
in_stream_full,
slice_stream_buff_0,
slice_stream_buff_1,
slice_stream_empty,
slice_stream_full,
stencil_stream_buff_0,
stencil_stream_buff_1,
stencil_stream_empty,
stencil_stream_full,
clk,rst,
step
);
input            arg_0_TREADY;
input      [7:0] arg_1_TDATA;
input            arg_1_TVALID;
input clk;
input rst;
input step;
output      [7:0] LB1D_buff;
output     [63:0] LB2D_proc_w;
output      [8:0] LB2D_proc_x;
output      [9:0] LB2D_proc_y;
output     [71:0] LB2D_shift_0;
output     [71:0] LB2D_shift_1;
output     [71:0] LB2D_shift_2;
output     [71:0] LB2D_shift_3;
output     [71:0] LB2D_shift_4;
output     [71:0] LB2D_shift_5;
output     [71:0] LB2D_shift_6;
output     [71:0] LB2D_shift_7;
output      [8:0] LB2D_shift_x;
output      [9:0] LB2D_shift_y;
output      [7:0] arg_0_TDATA;
output            arg_0_TVALID;
output            arg_1_TREADY;
output      [7:0] in_stream_buff_0;
output      [7:0] in_stream_buff_1;
output            in_stream_empty;
output            in_stream_full;
output     [71:0] slice_stream_buff_0;
output     [71:0] slice_stream_buff_1;
output            slice_stream_empty;
output            slice_stream_full;
output    [647:0] stencil_stream_buff_0;
output    [647:0] stencil_stream_buff_1;
output            stencil_stream_empty;
output            stencil_stream_full;
reg      [7:0] LB1D_buff;
reg     [63:0] LB2D_proc_w;
reg      [8:0] LB2D_proc_x;
reg      [9:0] LB2D_proc_y;
reg     [71:0] LB2D_shift_0;
reg     [71:0] LB2D_shift_1;
reg     [71:0] LB2D_shift_2;
reg     [71:0] LB2D_shift_3;
reg     [71:0] LB2D_shift_4;
reg     [71:0] LB2D_shift_5;
reg     [71:0] LB2D_shift_6;
reg     [71:0] LB2D_shift_7;
reg      [8:0] LB2D_shift_x;
reg      [9:0] LB2D_shift_y;
reg      [7:0] arg_0_TDATA;
reg            arg_0_TVALID;
reg            arg_1_TREADY;
reg      [7:0] in_stream_buff_0;
reg      [7:0] in_stream_buff_1;
reg            in_stream_empty;
reg            in_stream_full;
reg     [71:0] slice_stream_buff_0;
reg     [71:0] slice_stream_buff_1;
reg            slice_stream_empty;
reg            slice_stream_full;
reg    [647:0] stencil_stream_buff_0;
reg    [647:0] stencil_stream_buff_1;
reg            stencil_stream_empty;
reg            stencil_stream_full;
wire            arg_0_TREADY;
wire      [7:0] arg_1_TDATA;
wire            arg_1_TVALID;
wire            n0;
wire            n1;
wire            n2;
wire            n3;
wire            n4;
wire            n5;
wire            n6;
wire            n7;
wire            n8;
wire            n9;
wire            n10;
wire            n11;
wire            n12;
wire            n13;
wire            n14;
wire            n15;
wire      [7:0] n16;
wire      [7:0] n17;
wire      [7:0] n18;
wire      [7:0] n19;
wire            n20;
wire            n21;
wire     [63:0] n22;
wire     [63:0] n23;
wire     [63:0] n24;
wire     [63:0] n25;
wire     [63:0] n26;
wire     [63:0] n27;
wire     [63:0] n28;
wire      [8:0] n29;
wire      [8:0] n30;
wire      [8:0] n31;
wire      [8:0] n32;
wire      [8:0] n33;
wire      [8:0] n34;
wire            n35;
wire      [9:0] n36;
wire      [9:0] n37;
wire      [9:0] n38;
wire      [9:0] n39;
wire      [9:0] n40;
wire      [9:0] n41;
wire      [9:0] n42;
wire     [71:0] n43;
wire     [71:0] n44;
wire     [71:0] n45;
wire     [71:0] n46;
wire     [71:0] n47;
wire     [71:0] n48;
wire     [71:0] n49;
wire     [71:0] n50;
wire     [71:0] n51;
wire     [71:0] n52;
wire     [71:0] n53;
wire     [71:0] n54;
wire     [71:0] n55;
wire     [71:0] n56;
wire     [71:0] n57;
wire     [71:0] n58;
wire     [71:0] n59;
wire     [71:0] n60;
wire     [71:0] n61;
wire     [71:0] n62;
wire     [71:0] n63;
wire     [71:0] n64;
wire     [71:0] n65;
wire     [71:0] n66;
wire     [71:0] n67;
wire     [71:0] n68;
wire     [71:0] n69;
wire     [71:0] n70;
wire     [71:0] n71;
wire     [71:0] n72;
wire     [71:0] n73;
wire     [71:0] n74;
wire      [8:0] n75;
wire      [8:0] n76;
wire      [8:0] n77;
wire      [8:0] n78;
wire      [9:0] n79;
wire      [9:0] n80;
wire      [9:0] n81;
wire      [9:0] n82;
wire      [7:0] n83;
wire      [7:0] n84;
wire      [7:0] n85;
wire      [7:0] n86;
wire            n87;
wire            n88;
wire            n89;
wire            n90;
wire            n91;
wire            n92;
wire            n93;
wire            n94;
wire      [7:0] n95;
wire      [7:0] n96;
wire      [7:0] n97;
wire      [7:0] n98;
wire      [7:0] n99;
wire      [7:0] n100;
wire      [7:0] n101;
wire      [7:0] n102;
wire            n103;
wire            n104;
wire            n105;
wire            n106;
wire            n107;
wire            n108;
wire            n109;
wire            n110;
wire            n111;
wire            n112;
wire            n113;
wire            n114;
wire            n115;
wire      [7:0] n116;
wire            n117;
wire      [7:0] n118;
wire            n119;
wire      [7:0] n120;
wire            n121;
wire      [7:0] n122;
wire            n123;
wire      [7:0] n124;
wire            n125;
wire      [7:0] n126;
wire            n127;
wire      [7:0] n128;
wire            n129;
wire      [7:0] n130;
wire      [7:0] n131;
wire      [7:0] n132;
wire      [7:0] n133;
wire      [7:0] n134;
wire      [7:0] n135;
wire      [7:0] n136;
wire      [7:0] n137;
wire      [7:0] n138;
wire      [7:0] n139;
wire      [7:0] n140;
wire      [7:0] n141;
wire      [7:0] n142;
wire      [7:0] n143;
wire      [7:0] n144;
wire      [7:0] n145;
wire      [7:0] n146;
wire      [7:0] n147;
wire      [7:0] n148;
wire      [7:0] n149;
wire      [7:0] n150;
wire      [7:0] n151;
wire      [7:0] n152;
wire      [7:0] n153;
wire      [7:0] n154;
wire      [7:0] n155;
wire      [7:0] n156;
wire      [7:0] n157;
wire      [7:0] n158;
wire      [7:0] n159;
wire      [7:0] n160;
wire      [7:0] n161;
wire      [7:0] n162;
wire      [7:0] n163;
wire      [7:0] n164;
wire      [7:0] n165;
wire      [7:0] n166;
wire      [7:0] n167;
wire      [7:0] n168;
wire      [7:0] n169;
wire      [7:0] n170;
wire      [7:0] n171;
wire      [7:0] n172;
wire      [7:0] n173;
wire      [7:0] n174;
wire      [7:0] n175;
wire      [7:0] n176;
wire      [7:0] n177;
wire      [7:0] n178;
wire      [7:0] n179;
wire      [7:0] n180;
wire      [7:0] n181;
wire      [7:0] n182;
wire      [7:0] n183;
wire      [7:0] n184;
wire      [7:0] n185;
wire      [7:0] n186;
wire      [7:0] n187;
wire     [15:0] n188;
wire     [23:0] n189;
wire     [31:0] n190;
wire     [39:0] n191;
wire     [47:0] n192;
wire     [55:0] n193;
wire     [63:0] n194;
wire     [71:0] n195;
wire     [71:0] n196;
wire     [71:0] n197;
wire     [71:0] n198;
wire     [71:0] n199;
wire     [71:0] n200;
wire     [71:0] n201;
wire     [71:0] n202;
wire     [71:0] n203;
wire     [71:0] n204;
wire            n205;
wire            n206;
wire            n207;
wire            n208;
wire            n209;
wire            n210;
wire            n211;
wire            n212;
wire            n213;
wire            n214;
wire            n215;
wire            n216;
wire    [647:0] n217;
wire    [647:0] n218;
wire    [647:0] n219;
wire    [647:0] n220;
wire    [647:0] n221;
wire    [647:0] n222;
wire    [647:0] n223;
wire    [647:0] n224;
wire            n225;
wire            n226;
wire            n227;
wire            n228;
wire            n229;
wire            n230;
wire            n231;
wire            n232;
wire      [8:0] LB2D_proc_0_addr0;
wire      [7:0] LB2D_proc_0_data0;
wire            n233;
wire            n234;
wire            n235;
wire            n236;
wire            n237;
wire            n238;
wire            n239;
wire            n240;
wire            n241;
wire            n242;
wire            n243;
wire            n244;
wire            n245;
wire      [8:0] LB2D_proc_1_addr0;
wire      [7:0] LB2D_proc_1_data0;
wire            n246;
wire            n247;
wire            n248;
wire      [8:0] LB2D_proc_2_addr0;
wire      [7:0] LB2D_proc_2_data0;
wire            n249;
wire            n250;
wire            n251;
wire      [8:0] LB2D_proc_3_addr0;
wire      [7:0] LB2D_proc_3_data0;
wire            n252;
wire            n253;
wire            n254;
wire      [8:0] LB2D_proc_4_addr0;
wire      [7:0] LB2D_proc_4_data0;
wire            n255;
wire            n256;
wire            n257;
wire      [8:0] LB2D_proc_5_addr0;
wire      [7:0] LB2D_proc_5_data0;
wire            n258;
wire            n259;
wire            n260;
wire      [8:0] LB2D_proc_6_addr0;
wire      [7:0] LB2D_proc_6_data0;
wire            n261;
wire            n262;
wire            n263;
wire      [8:0] LB2D_proc_7_addr0;
wire      [7:0] LB2D_proc_7_data0;
wire            n264;
wire            n265;
wire            n266;
wire            n267;
reg      [7:0] LB2D_proc_0[511:0];
reg      [7:0] LB2D_proc_1[511:0];
reg      [7:0] LB2D_proc_2[511:0];
reg      [7:0] LB2D_proc_3[511:0];
reg      [7:0] LB2D_proc_4[511:0];
reg      [7:0] LB2D_proc_5[511:0];
reg      [7:0] LB2D_proc_6[511:0];
reg      [7:0] LB2D_proc_7[511:0];
wire clk;
wire rst;
wire step;
assign n0 =  ( in_stream_empty ) == ( 1'd0 )  ;
assign n1 =  ( slice_stream_full ) == ( 1'd0 )  ;
assign n2 =  ( n0 ) & ( n1 )  ;
assign n3 =  ( arg_1_TREADY ) == ( 1'd0 )  ;
assign n4 =  ( in_stream_full ) == ( 1'd0 )  ;
assign n5 =  ( n3 ) & ( n4 )  ;
assign n6 =  ( arg_0_TREADY ) == ( 1'd1 )  ;
assign n7 =  ( arg_0_TVALID ) == ( 1'd1 )  ;
assign n8 =  ( n6 ) & ( n7 )  ;
assign n9 =  ( arg_1_TVALID ) == ( 1'd0 )  ;
assign n10 =  ( n8 ) & ( n9 )  ;
assign n11 =  ( arg_1_TREADY ) == ( 1'd1 )  ;
assign n12 =  ( arg_1_TVALID ) == ( 1'd1 )  ;
assign n13 =  ( n11 ) & ( n12 )  ;
assign n14 =  ( arg_0_TREADY ) == ( 1'd0 )  ;
assign n15 =  ( n13 ) & ( n14 )  ;
assign n16 =  ( n15 ) ? ( arg_1_TDATA ) : ( LB1D_buff ) ;
assign n17 =  ( n10 ) ? ( arg_1_TDATA ) : ( n16 ) ;
assign n18 =  ( n5 ) ? ( LB1D_buff ) : ( n17 ) ;
assign n19 =  ( n2 ) ? ( LB1D_buff ) : ( n18 ) ;
assign n20 =  ( LB2D_proc_w ) < ( 64'd7 )  ;
assign n21 =  ( LB2D_proc_x ) < ( 9'd487 )  ;
assign n22 =  ( LB2D_proc_w ) + ( 64'd1 )  ;
assign n23 =  ( n21 ) ? ( LB2D_proc_w ) : ( n22 ) ;
assign n24 =  ( n20 ) ? ( n23 ) : ( 64'd0 ) ;
assign n25 =  ( n15 ) ? ( LB2D_proc_w ) : ( LB2D_proc_w ) ;
assign n26 =  ( n10 ) ? ( LB2D_proc_w ) : ( n25 ) ;
assign n27 =  ( n5 ) ? ( LB2D_proc_w ) : ( n26 ) ;
assign n28 =  ( n2 ) ? ( n24 ) : ( n27 ) ;
assign n29 =  ( LB2D_proc_x ) + ( 9'd1 )  ;
assign n30 =  ( n21 ) ? ( n29 ) : ( 9'd0 ) ;
assign n31 =  ( n15 ) ? ( LB2D_proc_x ) : ( LB2D_proc_x ) ;
assign n32 =  ( n10 ) ? ( LB2D_proc_x ) : ( n31 ) ;
assign n33 =  ( n5 ) ? ( LB2D_proc_x ) : ( n32 ) ;
assign n34 =  ( n2 ) ? ( n30 ) : ( n33 ) ;
assign n35 =  ( LB2D_proc_y ) < ( 10'd487 )  ;
assign n36 =  ( LB2D_proc_y ) + ( 10'd1 )  ;
assign n37 =  ( n21 ) ? ( LB2D_proc_y ) : ( n36 ) ;
assign n38 =  ( n35 ) ? ( n37 ) : ( 10'd487 ) ;
assign n39 =  ( n15 ) ? ( LB2D_proc_y ) : ( LB2D_proc_y ) ;
assign n40 =  ( n10 ) ? ( LB2D_proc_y ) : ( n39 ) ;
assign n41 =  ( n5 ) ? ( LB2D_proc_y ) : ( n40 ) ;
assign n42 =  ( n2 ) ? ( n38 ) : ( n41 ) ;
assign n43 =  ( n15 ) ? ( LB2D_shift_0 ) : ( LB2D_shift_0 ) ;
assign n44 =  ( n10 ) ? ( LB2D_shift_0 ) : ( n43 ) ;
assign n45 =  ( n5 ) ? ( LB2D_shift_0 ) : ( n44 ) ;
assign n46 =  ( n2 ) ? ( LB2D_shift_0 ) : ( n45 ) ;
assign n47 =  ( n15 ) ? ( LB2D_shift_1 ) : ( LB2D_shift_1 ) ;
assign n48 =  ( n10 ) ? ( LB2D_shift_1 ) : ( n47 ) ;
assign n49 =  ( n5 ) ? ( LB2D_shift_1 ) : ( n48 ) ;
assign n50 =  ( n2 ) ? ( LB2D_shift_1 ) : ( n49 ) ;
assign n51 =  ( n15 ) ? ( LB2D_shift_2 ) : ( LB2D_shift_2 ) ;
assign n52 =  ( n10 ) ? ( LB2D_shift_2 ) : ( n51 ) ;
assign n53 =  ( n5 ) ? ( LB2D_shift_2 ) : ( n52 ) ;
assign n54 =  ( n2 ) ? ( LB2D_shift_2 ) : ( n53 ) ;
assign n55 =  ( n15 ) ? ( LB2D_shift_3 ) : ( LB2D_shift_3 ) ;
assign n56 =  ( n10 ) ? ( LB2D_shift_3 ) : ( n55 ) ;
assign n57 =  ( n5 ) ? ( LB2D_shift_3 ) : ( n56 ) ;
assign n58 =  ( n2 ) ? ( LB2D_shift_3 ) : ( n57 ) ;
assign n59 =  ( n15 ) ? ( LB2D_shift_4 ) : ( LB2D_shift_4 ) ;
assign n60 =  ( n10 ) ? ( LB2D_shift_4 ) : ( n59 ) ;
assign n61 =  ( n5 ) ? ( LB2D_shift_4 ) : ( n60 ) ;
assign n62 =  ( n2 ) ? ( LB2D_shift_4 ) : ( n61 ) ;
assign n63 =  ( n15 ) ? ( LB2D_shift_5 ) : ( LB2D_shift_5 ) ;
assign n64 =  ( n10 ) ? ( LB2D_shift_5 ) : ( n63 ) ;
assign n65 =  ( n5 ) ? ( LB2D_shift_5 ) : ( n64 ) ;
assign n66 =  ( n2 ) ? ( LB2D_shift_5 ) : ( n65 ) ;
assign n67 =  ( n15 ) ? ( LB2D_shift_6 ) : ( LB2D_shift_6 ) ;
assign n68 =  ( n10 ) ? ( LB2D_shift_6 ) : ( n67 ) ;
assign n69 =  ( n5 ) ? ( LB2D_shift_6 ) : ( n68 ) ;
assign n70 =  ( n2 ) ? ( LB2D_shift_6 ) : ( n69 ) ;
assign n71 =  ( n15 ) ? ( LB2D_shift_7 ) : ( LB2D_shift_7 ) ;
assign n72 =  ( n10 ) ? ( LB2D_shift_7 ) : ( n71 ) ;
assign n73 =  ( n5 ) ? ( LB2D_shift_7 ) : ( n72 ) ;
assign n74 =  ( n2 ) ? ( LB2D_shift_7 ) : ( n73 ) ;
assign n75 =  ( n15 ) ? ( LB2D_shift_x ) : ( LB2D_shift_x ) ;
assign n76 =  ( n10 ) ? ( LB2D_shift_x ) : ( n75 ) ;
assign n77 =  ( n5 ) ? ( LB2D_shift_x ) : ( n76 ) ;
assign n78 =  ( n2 ) ? ( LB2D_shift_x ) : ( n77 ) ;
assign n79 =  ( n15 ) ? ( LB2D_shift_y ) : ( LB2D_shift_y ) ;
assign n80 =  ( n10 ) ? ( LB2D_shift_y ) : ( n79 ) ;
assign n81 =  ( n5 ) ? ( LB2D_shift_y ) : ( n80 ) ;
assign n82 =  ( n2 ) ? ( LB2D_shift_y ) : ( n81 ) ;
assign n83 =  ( n15 ) ? ( arg_0_TDATA ) : ( arg_0_TDATA ) ;
assign n84 =  ( n10 ) ? ( arg_0_TDATA ) : ( n83 ) ;
assign n85 =  ( n5 ) ? ( arg_0_TDATA ) : ( n84 ) ;
assign n86 =  ( n2 ) ? ( arg_0_TDATA ) : ( n85 ) ;
assign n87 =  ( n15 ) ? ( arg_0_TVALID ) : ( arg_0_TVALID ) ;
assign n88 =  ( n10 ) ? ( 1'd0 ) : ( n87 ) ;
assign n89 =  ( n5 ) ? ( arg_0_TVALID ) : ( n88 ) ;
assign n90 =  ( n2 ) ? ( arg_0_TVALID ) : ( n89 ) ;
assign n91 =  ( n15 ) ? ( 1'd0 ) : ( arg_1_TREADY ) ;
assign n92 =  ( n10 ) ? ( 1'd0 ) : ( n91 ) ;
assign n93 =  ( n5 ) ? ( 1'd1 ) : ( n92 ) ;
assign n94 =  ( n2 ) ? ( arg_1_TREADY ) : ( n93 ) ;
assign n95 =  ( n15 ) ? ( in_stream_buff_0 ) : ( in_stream_buff_0 ) ;
assign n96 =  ( n10 ) ? ( in_stream_buff_0 ) : ( n95 ) ;
assign n97 =  ( n5 ) ? ( LB1D_buff ) : ( n96 ) ;
assign n98 =  ( n2 ) ? ( in_stream_buff_0 ) : ( n97 ) ;
assign n99 =  ( n15 ) ? ( in_stream_buff_1 ) : ( in_stream_buff_1 ) ;
assign n100 =  ( n10 ) ? ( in_stream_buff_1 ) : ( n99 ) ;
assign n101 =  ( n5 ) ? ( in_stream_buff_0 ) : ( n100 ) ;
assign n102 =  ( n2 ) ? ( in_stream_buff_1 ) : ( n101 ) ;
assign n103 =  ( in_stream_full ) == ( 1'd1 )  ;
assign n104 =  ( n103 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n105 =  ( n15 ) ? ( in_stream_empty ) : ( in_stream_empty ) ;
assign n106 =  ( n10 ) ? ( in_stream_empty ) : ( n105 ) ;
assign n107 =  ( n5 ) ? ( 1'd0 ) : ( n106 ) ;
assign n108 =  ( n2 ) ? ( n104 ) : ( n107 ) ;
assign n109 =  ( in_stream_empty ) == ( 1'd1 )  ;
assign n110 =  ( n109 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n111 =  ( n15 ) ? ( in_stream_full ) : ( in_stream_full ) ;
assign n112 =  ( n10 ) ? ( in_stream_full ) : ( n111 ) ;
assign n113 =  ( n5 ) ? ( n110 ) : ( n112 ) ;
assign n114 =  ( n2 ) ? ( 1'd0 ) : ( n113 ) ;
assign n115 =  ( LB2D_proc_y ) >= ( 10'd8 )  ;
assign n116 =  ( n103 ) ? ( in_stream_buff_1 ) : ( in_stream_buff_0 ) ;
assign n117 =  ( LB2D_proc_w ) == ( 64'd0 )  ;
assign n118 =  (  LB2D_proc_7 [ LB2D_proc_x ] )  ;
assign n119 =  ( LB2D_proc_w ) == ( 64'd1 )  ;
assign n120 =  (  LB2D_proc_0 [ LB2D_proc_x ] )  ;
assign n121 =  ( LB2D_proc_w ) == ( 64'd2 )  ;
assign n122 =  (  LB2D_proc_1 [ LB2D_proc_x ] )  ;
assign n123 =  ( LB2D_proc_w ) == ( 64'd3 )  ;
assign n124 =  (  LB2D_proc_2 [ LB2D_proc_x ] )  ;
assign n125 =  ( LB2D_proc_w ) == ( 64'd4 )  ;
assign n126 =  (  LB2D_proc_3 [ LB2D_proc_x ] )  ;
assign n127 =  ( LB2D_proc_w ) == ( 64'd5 )  ;
assign n128 =  (  LB2D_proc_4 [ LB2D_proc_x ] )  ;
assign n129 =  ( LB2D_proc_w ) == ( 64'd6 )  ;
assign n130 =  (  LB2D_proc_5 [ LB2D_proc_x ] )  ;
assign n131 =  (  LB2D_proc_6 [ LB2D_proc_x ] )  ;
assign n132 =  ( n129 ) ? ( n130 ) : ( n131 ) ;
assign n133 =  ( n127 ) ? ( n128 ) : ( n132 ) ;
assign n134 =  ( n125 ) ? ( n126 ) : ( n133 ) ;
assign n135 =  ( n123 ) ? ( n124 ) : ( n134 ) ;
assign n136 =  ( n121 ) ? ( n122 ) : ( n135 ) ;
assign n137 =  ( n119 ) ? ( n120 ) : ( n136 ) ;
assign n138 =  ( n117 ) ? ( n118 ) : ( n137 ) ;
assign n139 =  ( n129 ) ? ( n128 ) : ( n130 ) ;
assign n140 =  ( n127 ) ? ( n126 ) : ( n139 ) ;
assign n141 =  ( n125 ) ? ( n124 ) : ( n140 ) ;
assign n142 =  ( n123 ) ? ( n122 ) : ( n141 ) ;
assign n143 =  ( n121 ) ? ( n120 ) : ( n142 ) ;
assign n144 =  ( n119 ) ? ( n118 ) : ( n143 ) ;
assign n145 =  ( n117 ) ? ( n131 ) : ( n144 ) ;
assign n146 =  ( n129 ) ? ( n126 ) : ( n128 ) ;
assign n147 =  ( n127 ) ? ( n124 ) : ( n146 ) ;
assign n148 =  ( n125 ) ? ( n122 ) : ( n147 ) ;
assign n149 =  ( n123 ) ? ( n120 ) : ( n148 ) ;
assign n150 =  ( n121 ) ? ( n118 ) : ( n149 ) ;
assign n151 =  ( n119 ) ? ( n131 ) : ( n150 ) ;
assign n152 =  ( n117 ) ? ( n130 ) : ( n151 ) ;
assign n153 =  ( n129 ) ? ( n124 ) : ( n126 ) ;
assign n154 =  ( n127 ) ? ( n122 ) : ( n153 ) ;
assign n155 =  ( n125 ) ? ( n120 ) : ( n154 ) ;
assign n156 =  ( n123 ) ? ( n118 ) : ( n155 ) ;
assign n157 =  ( n121 ) ? ( n131 ) : ( n156 ) ;
assign n158 =  ( n119 ) ? ( n130 ) : ( n157 ) ;
assign n159 =  ( n117 ) ? ( n128 ) : ( n158 ) ;
assign n160 =  ( n129 ) ? ( n122 ) : ( n124 ) ;
assign n161 =  ( n127 ) ? ( n120 ) : ( n160 ) ;
assign n162 =  ( n125 ) ? ( n118 ) : ( n161 ) ;
assign n163 =  ( n123 ) ? ( n131 ) : ( n162 ) ;
assign n164 =  ( n121 ) ? ( n130 ) : ( n163 ) ;
assign n165 =  ( n119 ) ? ( n128 ) : ( n164 ) ;
assign n166 =  ( n117 ) ? ( n126 ) : ( n165 ) ;
assign n167 =  ( n129 ) ? ( n120 ) : ( n122 ) ;
assign n168 =  ( n127 ) ? ( n118 ) : ( n167 ) ;
assign n169 =  ( n125 ) ? ( n131 ) : ( n168 ) ;
assign n170 =  ( n123 ) ? ( n130 ) : ( n169 ) ;
assign n171 =  ( n121 ) ? ( n128 ) : ( n170 ) ;
assign n172 =  ( n119 ) ? ( n126 ) : ( n171 ) ;
assign n173 =  ( n117 ) ? ( n124 ) : ( n172 ) ;
assign n174 =  ( n129 ) ? ( n118 ) : ( n120 ) ;
assign n175 =  ( n127 ) ? ( n131 ) : ( n174 ) ;
assign n176 =  ( n125 ) ? ( n130 ) : ( n175 ) ;
assign n177 =  ( n123 ) ? ( n128 ) : ( n176 ) ;
assign n178 =  ( n121 ) ? ( n126 ) : ( n177 ) ;
assign n179 =  ( n119 ) ? ( n124 ) : ( n178 ) ;
assign n180 =  ( n117 ) ? ( n122 ) : ( n179 ) ;
assign n181 =  ( n129 ) ? ( n131 ) : ( n118 ) ;
assign n182 =  ( n127 ) ? ( n130 ) : ( n181 ) ;
assign n183 =  ( n125 ) ? ( n128 ) : ( n182 ) ;
assign n184 =  ( n123 ) ? ( n126 ) : ( n183 ) ;
assign n185 =  ( n121 ) ? ( n124 ) : ( n184 ) ;
assign n186 =  ( n119 ) ? ( n122 ) : ( n185 ) ;
assign n187 =  ( n117 ) ? ( n120 ) : ( n186 ) ;
assign n188 =  { ( n180 ) , ( n187 ) }  ;
assign n189 =  { ( n173 ) , ( n188 ) }  ;
assign n190 =  { ( n166 ) , ( n189 ) }  ;
assign n191 =  { ( n159 ) , ( n190 ) }  ;
assign n192 =  { ( n152 ) , ( n191 ) }  ;
assign n193 =  { ( n145 ) , ( n192 ) }  ;
assign n194 =  { ( n138 ) , ( n193 ) }  ;
assign n195 =  { ( n116 ) , ( n194 ) }  ;
assign n196 =  ( n115 ) ? ( n195 ) : ( slice_stream_buff_0 ) ;
assign n197 =  ( n15 ) ? ( slice_stream_buff_0 ) : ( slice_stream_buff_0 ) ;
assign n198 =  ( n10 ) ? ( slice_stream_buff_0 ) : ( n197 ) ;
assign n199 =  ( n5 ) ? ( slice_stream_buff_0 ) : ( n198 ) ;
assign n200 =  ( n2 ) ? ( n196 ) : ( n199 ) ;
assign n201 =  ( n15 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_1 ) ;
assign n202 =  ( n10 ) ? ( slice_stream_buff_1 ) : ( n201 ) ;
assign n203 =  ( n5 ) ? ( slice_stream_buff_1 ) : ( n202 ) ;
assign n204 =  ( n2 ) ? ( slice_stream_buff_0 ) : ( n203 ) ;
assign n205 =  ( n115 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n206 =  ( n15 ) ? ( slice_stream_empty ) : ( slice_stream_empty ) ;
assign n207 =  ( n10 ) ? ( slice_stream_empty ) : ( n206 ) ;
assign n208 =  ( n5 ) ? ( slice_stream_empty ) : ( n207 ) ;
assign n209 =  ( n2 ) ? ( n205 ) : ( n208 ) ;
assign n210 =  ( slice_stream_empty ) == ( 1'd1 )  ;
assign n211 =  ( n210 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n212 =  ( n115 ) ? ( n211 ) : ( 1'd0 ) ;
assign n213 =  ( n15 ) ? ( slice_stream_full ) : ( slice_stream_full ) ;
assign n214 =  ( n10 ) ? ( slice_stream_full ) : ( n213 ) ;
assign n215 =  ( n5 ) ? ( slice_stream_full ) : ( n214 ) ;
assign n216 =  ( n2 ) ? ( n212 ) : ( n215 ) ;
assign n217 =  ( n15 ) ? ( stencil_stream_buff_0 ) : ( stencil_stream_buff_0 ) ;
assign n218 =  ( n10 ) ? ( stencil_stream_buff_0 ) : ( n217 ) ;
assign n219 =  ( n5 ) ? ( stencil_stream_buff_0 ) : ( n218 ) ;
assign n220 =  ( n2 ) ? ( stencil_stream_buff_0 ) : ( n219 ) ;
assign n221 =  ( n15 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_1 ) ;
assign n222 =  ( n10 ) ? ( stencil_stream_buff_1 ) : ( n221 ) ;
assign n223 =  ( n5 ) ? ( stencil_stream_buff_1 ) : ( n222 ) ;
assign n224 =  ( n2 ) ? ( stencil_stream_buff_1 ) : ( n223 ) ;
assign n225 =  ( n15 ) ? ( stencil_stream_empty ) : ( stencil_stream_empty ) ;
assign n226 =  ( n10 ) ? ( stencil_stream_empty ) : ( n225 ) ;
assign n227 =  ( n5 ) ? ( stencil_stream_empty ) : ( n226 ) ;
assign n228 =  ( n2 ) ? ( stencil_stream_empty ) : ( n227 ) ;
assign n229 =  ( n15 ) ? ( stencil_stream_full ) : ( stencil_stream_full ) ;
assign n230 =  ( n10 ) ? ( stencil_stream_full ) : ( n229 ) ;
assign n231 =  ( n5 ) ? ( stencil_stream_full ) : ( n230 ) ;
assign n232 =  ( n2 ) ? ( stencil_stream_full ) : ( n231 ) ;
assign n233 = ~ ( n2 ) ;
assign n234 = ~ ( n5 ) ;
assign n235 =  ( n233 ) & ( n234 )  ;
assign n236 = ~ ( n10 ) ;
assign n237 =  ( n235 ) & ( n236 )  ;
assign n238 = ~ ( n15 ) ;
assign n239 =  ( n237 ) & ( n238 )  ;
assign n240 =  ( n237 ) & ( n15 )  ;
assign n241 =  ( n235 ) & ( n10 )  ;
assign n242 =  ( n233 ) & ( n5 )  ;
assign n243 = ~ ( n117 ) ;
assign n244 =  ( n2 ) & ( n243 )  ;
assign n245 =  ( n2 ) & ( n117 )  ;
assign LB2D_proc_0_addr0 = n245 ? (LB2D_proc_x) : (0);
assign LB2D_proc_0_data0 = n245 ? (n116) : (LB2D_proc_0[0]);
assign n246 = ~ ( n119 ) ;
assign n247 =  ( n2 ) & ( n246 )  ;
assign n248 =  ( n2 ) & ( n119 )  ;
assign LB2D_proc_1_addr0 = n248 ? (LB2D_proc_x) : (0);
assign LB2D_proc_1_data0 = n248 ? (n116) : (LB2D_proc_1[0]);
assign n249 = ~ ( n121 ) ;
assign n250 =  ( n2 ) & ( n249 )  ;
assign n251 =  ( n2 ) & ( n121 )  ;
assign LB2D_proc_2_addr0 = n251 ? (LB2D_proc_x) : (0);
assign LB2D_proc_2_data0 = n251 ? (n116) : (LB2D_proc_2[0]);
assign n252 = ~ ( n123 ) ;
assign n253 =  ( n2 ) & ( n252 )  ;
assign n254 =  ( n2 ) & ( n123 )  ;
assign LB2D_proc_3_addr0 = n254 ? (LB2D_proc_x) : (0);
assign LB2D_proc_3_data0 = n254 ? (n116) : (LB2D_proc_3[0]);
assign n255 = ~ ( n125 ) ;
assign n256 =  ( n2 ) & ( n255 )  ;
assign n257 =  ( n2 ) & ( n125 )  ;
assign LB2D_proc_4_addr0 = n257 ? (LB2D_proc_x) : (0);
assign LB2D_proc_4_data0 = n257 ? (n116) : (LB2D_proc_4[0]);
assign n258 = ~ ( n127 ) ;
assign n259 =  ( n2 ) & ( n258 )  ;
assign n260 =  ( n2 ) & ( n127 )  ;
assign LB2D_proc_5_addr0 = n260 ? (LB2D_proc_x) : (0);
assign LB2D_proc_5_data0 = n260 ? (n116) : (LB2D_proc_5[0]);
assign n261 = ~ ( n129 ) ;
assign n262 =  ( n2 ) & ( n261 )  ;
assign n263 =  ( n2 ) & ( n129 )  ;
assign LB2D_proc_6_addr0 = n263 ? (LB2D_proc_x) : (0);
assign LB2D_proc_6_data0 = n263 ? (n116) : (LB2D_proc_6[0]);
assign n264 =  ( LB2D_proc_w ) == ( 64'd7 )  ;
assign n265 = ~ ( n264 ) ;
assign n266 =  ( n2 ) & ( n265 )  ;
assign n267 =  ( n2 ) & ( n264 )  ;
assign LB2D_proc_7_addr0 = n267 ? (LB2D_proc_x) : (0);
assign LB2D_proc_7_data0 = n267 ? (n116) : (LB2D_proc_7[0]);
always @(posedge clk) begin
   if(rst) begin
       LB1D_buff <= LB1D_buff;
       LB2D_proc_w <= LB2D_proc_w;
       LB2D_proc_x <= LB2D_proc_x;
       LB2D_proc_y <= LB2D_proc_y;
       LB2D_shift_0 <= LB2D_shift_0;
       LB2D_shift_1 <= LB2D_shift_1;
       LB2D_shift_2 <= LB2D_shift_2;
       LB2D_shift_3 <= LB2D_shift_3;
       LB2D_shift_4 <= LB2D_shift_4;
       LB2D_shift_5 <= LB2D_shift_5;
       LB2D_shift_6 <= LB2D_shift_6;
       LB2D_shift_7 <= LB2D_shift_7;
       LB2D_shift_x <= LB2D_shift_x;
       LB2D_shift_y <= LB2D_shift_y;
       arg_0_TDATA <= arg_0_TDATA;
       arg_0_TVALID <= arg_0_TVALID;
       arg_1_TREADY <= arg_1_TREADY;
       in_stream_buff_0 <= in_stream_buff_0;
       in_stream_buff_1 <= in_stream_buff_1;
       in_stream_empty <= in_stream_empty;
       in_stream_full <= in_stream_full;
       slice_stream_buff_0 <= slice_stream_buff_0;
       slice_stream_buff_1 <= slice_stream_buff_1;
       slice_stream_empty <= slice_stream_empty;
       slice_stream_full <= slice_stream_full;
       stencil_stream_buff_0 <= stencil_stream_buff_0;
       stencil_stream_buff_1 <= stencil_stream_buff_1;
       stencil_stream_empty <= stencil_stream_empty;
       stencil_stream_full <= stencil_stream_full;
   end
   else if(step) begin
       LB1D_buff <= n19;
       LB2D_proc_w <= n28;
       LB2D_proc_x <= n34;
       LB2D_proc_y <= n42;
       LB2D_shift_0 <= n46;
       LB2D_shift_1 <= n50;
       LB2D_shift_2 <= n54;
       LB2D_shift_3 <= n58;
       LB2D_shift_4 <= n62;
       LB2D_shift_5 <= n66;
       LB2D_shift_6 <= n70;
       LB2D_shift_7 <= n74;
       LB2D_shift_x <= n78;
       LB2D_shift_y <= n82;
       arg_0_TDATA <= n86;
       arg_0_TVALID <= n90;
       arg_1_TREADY <= n94;
       in_stream_buff_0 <= n98;
       in_stream_buff_1 <= n102;
       in_stream_empty <= n108;
       in_stream_full <= n114;
       slice_stream_buff_0 <= n200;
       slice_stream_buff_1 <= n204;
       slice_stream_empty <= n209;
       slice_stream_full <= n216;
       stencil_stream_buff_0 <= n220;
       stencil_stream_buff_1 <= n224;
       stencil_stream_empty <= n228;
       stencil_stream_full <= n232;
       LB2D_proc_0 [ LB2D_proc_0_addr0 ] <= LB2D_proc_0_data0;
       LB2D_proc_1 [ LB2D_proc_1_addr0 ] <= LB2D_proc_1_data0;
       LB2D_proc_2 [ LB2D_proc_2_addr0 ] <= LB2D_proc_2_data0;
       LB2D_proc_3 [ LB2D_proc_3_addr0 ] <= LB2D_proc_3_data0;
       LB2D_proc_4 [ LB2D_proc_4_addr0 ] <= LB2D_proc_4_data0;
       LB2D_proc_5 [ LB2D_proc_5_addr0 ] <= LB2D_proc_5_data0;
       LB2D_proc_6 [ LB2D_proc_6_addr0 ] <= LB2D_proc_6_data0;
       LB2D_proc_7 [ LB2D_proc_7_addr0 ] <= LB2D_proc_7_data0;
   end
end
endmodule
