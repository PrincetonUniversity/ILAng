module riscv(
meInt,
msInt,
mtInt,
seInt,
ssInt,
stInt,
mem_data_n112,
mem_data_n1080,
mem_data_n2862,
Priv,
mbadaddr,
mcause,
medeleg,
mepc,
mideleg,
mie,
mip,
misa,
mscratch,
mstatus,
mtvec,
pc,
sbadaddr,
scause,
sepc,
sptbr,
sscratch,
stvec,
x0,
x1,
x10,
x11,
x12,
x13,
x14,
x15,
x16,
x17,
x18,
x19,
x2,
x20,
x21,
x22,
x23,
x24,
x25,
x26,
x27,
x28,
x29,
x3,
x30,
x31,
x4,
x5,
x6,
x7,
x8,
x9,
mem_addr_n111,
mem_addr_n1079,
mem_addr0,
mem_data0,
mem_wen0,
mem_addr_n2861,
clk,rst,
step
);
input            meInt;
input            msInt;
input            mtInt;
input            seInt;
input            ssInt;
input            stInt;
input     [31:0] mem_data_n112;
input     [31:0] mem_data_n1080;
input     [31:0] mem_data_n2862;
input clk;
input rst;
input step;
output      [1:0] Priv;
output     [31:0] mbadaddr;
output     [31:0] mcause;
output     [31:0] medeleg;
output     [31:0] mepc;
output     [31:0] mideleg;
output     [31:0] mie;
output     [31:0] mip;
output     [31:0] misa;
output     [31:0] mscratch;
output     [31:0] mstatus;
output     [31:0] mtvec;
output     [31:0] pc;
output     [31:0] sbadaddr;
output     [31:0] scause;
output     [31:0] sepc;
output     [31:0] sptbr;
output     [31:0] sscratch;
output     [31:0] stvec;
output     [31:0] x0;
output     [31:0] x1;
output     [31:0] x10;
output     [31:0] x11;
output     [31:0] x12;
output     [31:0] x13;
output     [31:0] x14;
output     [31:0] x15;
output     [31:0] x16;
output     [31:0] x17;
output     [31:0] x18;
output     [31:0] x19;
output     [31:0] x2;
output     [31:0] x20;
output     [31:0] x21;
output     [31:0] x22;
output     [31:0] x23;
output     [31:0] x24;
output     [31:0] x25;
output     [31:0] x26;
output     [31:0] x27;
output     [31:0] x28;
output     [31:0] x29;
output     [31:0] x3;
output     [31:0] x30;
output     [31:0] x31;
output     [31:0] x4;
output     [31:0] x5;
output     [31:0] x6;
output     [31:0] x7;
output     [31:0] x8;
output     [31:0] x9;
output     [31:0] mem_addr_n111;
output     [31:0] mem_addr_n1079;
output     [31:0] mem_addr0;
output     [31:0] mem_data0;
output            mem_wen0;
output     [31:0] mem_addr_n2861;
reg      [1:0] Priv;
reg     [31:0] mbadaddr;
reg     [31:0] mcause;
reg     [31:0] medeleg;
reg     [31:0] mepc;
reg     [31:0] mideleg;
reg     [31:0] mie;
reg     [31:0] mip;
reg     [31:0] misa;
reg     [31:0] mscratch;
reg     [31:0] mstatus;
reg     [31:0] mtvec;
reg     [31:0] pc;
reg     [31:0] sbadaddr;
reg     [31:0] scause;
reg     [31:0] sepc;
reg     [31:0] sptbr;
reg     [31:0] sscratch;
reg     [31:0] stvec;
reg     [31:0] x0;
reg     [31:0] x1;
reg     [31:0] x10;
reg     [31:0] x11;
reg     [31:0] x12;
reg     [31:0] x13;
reg     [31:0] x14;
reg     [31:0] x15;
reg     [31:0] x16;
reg     [31:0] x17;
reg     [31:0] x18;
reg     [31:0] x19;
reg     [31:0] x2;
reg     [31:0] x20;
reg     [31:0] x21;
reg     [31:0] x22;
reg     [31:0] x23;
reg     [31:0] x24;
reg     [31:0] x25;
reg     [31:0] x26;
reg     [31:0] x27;
reg     [31:0] x28;
reg     [31:0] x29;
reg     [31:0] x3;
reg     [31:0] x30;
reg     [31:0] x31;
reg     [31:0] x4;
reg     [31:0] x5;
reg     [31:0] x6;
reg     [31:0] x7;
reg     [31:0] x8;
reg     [31:0] x9;
wire            meInt;
wire            msInt;
wire            mtInt;
wire            seInt;
wire            ssInt;
wire            stInt;
wire            n0;
wire            n1;
wire            n2;
wire            n3;
wire            n4;
wire            n5;
wire      [1:0] n6;
wire      [2:0] n7;
wire      [3:0] n8;
wire      [4:0] n9;
wire      [5:0] n10;
wire      [6:0] n11;
wire      [7:0] n12;
wire      [8:0] n13;
wire      [9:0] n14;
wire     [10:0] n15;
wire     [11:0] n16;
wire     [31:0] n17;
wire     [31:0] n18;
wire            n19;
wire            n20;
wire            n21;
wire            n22;
wire            n23;
wire     [31:0] n24;
wire            n25;
wire            n26;
wire            n27;
wire            n28;
wire            n29;
wire            n30;
wire            n31;
wire            n32;
wire            n33;
wire            n34;
wire            n35;
wire            n36;
wire            n37;
wire            n38;
wire            n39;
wire            n40;
wire     [31:0] n41;
wire            n42;
wire            n43;
wire            n44;
wire            n45;
wire            n46;
wire     [31:0] n47;
wire            n48;
wire            n49;
wire            n50;
wire            n51;
wire            n52;
wire            n53;
wire            n54;
wire            n55;
wire            n56;
wire            n57;
wire     [31:0] n58;
wire            n59;
wire            n60;
wire            n61;
wire            n62;
wire            n63;
wire     [31:0] n64;
wire            n65;
wire            n66;
wire            n67;
wire            n68;
wire            n69;
wire            n70;
wire            n71;
wire            n72;
wire            n73;
wire            n74;
wire     [31:0] n75;
wire     [31:0] n76;
wire     [31:0] n77;
wire     [31:0] n78;
wire     [31:0] n79;
wire     [31:0] n80;
wire     [31:0] n81;
wire     [31:0] n82;
wire     [31:0] n83;
wire     [31:0] n84__int_trap_select;
wire            n85;
wire            n86;
wire            n87;
wire            n88;
wire            n89;
wire            n90;
wire            n91;
wire            n92;
wire            n93;
wire            n94;
wire            n95;
wire            n96;
wire            n97;
wire            n98;
wire            n99;
wire            n100;
wire            n101;
wire            n102;
wire            n103;
wire            n104;
wire            n105;
wire            n106__take_int_sig;
wire      [1:0] n107;
wire            n108;
wire     [29:0] n109;
wire     [31:0] n110;
wire     [31:0] n113;
wire            n114;
wire            n115;
wire            n116;
wire      [1:0] n117;
wire            n118;
wire            n119;
wire      [1:0] n120;
wire            n121;
wire            n122;
wire            n123;
wire            n124;
wire            n125;
wire     [31:0] n126;
wire            n127;
wire            n128;
wire            n129;
wire     [31:0] n130;
wire            n131;
wire            n132;
wire            n133;
wire            n134;
wire            n135;
wire            n136;
wire            n137;
wire            n138;
wire            n139;
wire     [31:0] n140;
wire            n141;
wire            n142;
wire            n143;
wire            n144;
wire            n145;
wire            n146;
wire     [31:0] n147;
wire            n148;
wire            n149;
wire            n150;
wire            n151;
wire            n152;
wire            n153;
wire            n154;
wire            n155;
wire            n156;
wire            n157;
wire            n158;
wire            n159;
wire            n160;
wire            n161;
wire     [31:0] n162;
wire            n163;
wire     [31:0] n164;
wire            n165;
wire            n166;
wire     [31:0] n167;
wire            n168;
wire            n169;
wire     [31:0] n170;
wire            n171;
wire            n172;
wire            n173;
wire            n174;
wire            n175;
wire            n176;
wire            n177;
wire            n178;
wire     [31:0] n179;
wire            n180;
wire            n181;
wire            n182;
wire            n183;
wire     [31:0] n184;
wire            n185;
wire     [31:0] n186;
wire            n187;
wire            n188;
wire            n189;
wire            n190;
wire            n191;
wire            n192;
wire            n193;
wire            n194;
wire            n195;
wire            n196;
wire            n197;
wire            n198;
wire            n199;
wire            n200;
wire            n201;
wire            n202;
wire            n203;
wire            n204;
wire            n205;
wire            n206;
wire            n207;
wire     [31:0] n208;
wire            n209;
wire            n210;
wire            n211;
wire            n212;
wire            n213;
wire            n214;
wire            n215;
wire            n216;
wire            n217;
wire            n218;
wire            n219;
wire            n220;
wire            n221;
wire            n222;
wire     [31:0] n223;
wire            n224;
wire            n225;
wire            n226;
wire            n227;
wire            n228;
wire            n229;
wire            n230;
wire            n231;
wire            n232;
wire            n233;
wire            n234;
wire            n235;
wire            n236;
wire            n237;
wire            n238;
wire            n239;
wire            n240;
wire            n241;
wire            n242;
wire            n243;
wire     [31:0] n244;
wire            n245;
wire     [31:0] n246;
wire            n247;
wire            n248;
wire            n249;
wire            n250;
wire            n251;
wire            n252;
wire            n253;
wire            n254;
wire     [31:0] n255;
wire            n256;
wire     [31:0] n257;
wire            n258;
wire            n259;
wire            n260;
wire            n261;
wire            n262;
wire            n263;
wire            n264;
wire            n265;
wire            n266;
wire            n267;
wire            n268;
wire            n269;
wire            n270;
wire            n271;
wire            n272;
wire            n273;
wire            n274;
wire            n275;
wire            n276;
wire            n277;
wire            n278;
wire            n279;
wire            n280;
wire            n281;
wire            n282;
wire            n283;
wire            n284;
wire            n285;
wire            n286;
wire            n287;
wire            n288;
wire            n289;
wire            n290;
wire            n291;
wire            n292;
wire            n293;
wire            n294;
wire            n295;
wire            n296;
wire            n297;
wire            n298;
wire            n299;
wire            n300;
wire            n301;
wire            n302;
wire            n303;
wire            n304;
wire            n305;
wire            n306;
wire            n307;
wire            n308;
wire            n309;
wire            n310;
wire            n311;
wire            n312;
wire            n313;
wire            n314;
wire            n315;
wire            n316;
wire            n317;
wire            n318;
wire            n319;
wire            n320;
wire            n321;
wire            n322;
wire            n323;
wire            n324;
wire            n325;
wire     [31:0] n326;
wire            n327;
wire            n328;
wire            n329;
wire            n330;
wire            n331;
wire            n332;
wire            n333;
wire     [31:0] n334;
wire            n335;
wire            n336;
wire            n337;
wire            n338;
wire            n339;
wire            n340;
wire            n341;
wire            n342;
wire            n343;
wire            n344;
wire            n345;
wire            n346;
wire            n347;
wire            n348;
wire            n349;
wire            n350;
wire            n351;
wire            n352;
wire            n353;
wire            n354;
wire            n355;
wire            n356;
wire            n357;
wire            n358;
wire            n359;
wire            n360;
wire            n361;
wire            n362;
wire            n363;
wire            n364;
wire            n365;
wire            n366;
wire            n367;
wire            n368;
wire            n369;
wire            n370;
wire            n371;
wire            n372;
wire            n373;
wire            n374;
wire            n375;
wire            n376;
wire            n377;
wire            n378;
wire            n379;
wire            n380;
wire            n381;
wire            n382;
wire            n383;
wire            n384;
wire            n385;
wire            n386;
wire            n387;
wire            n388;
wire            n389;
wire            n390;
wire            n391;
wire            n392;
wire            n393;
wire            n394;
wire            n395;
wire            n396;
wire            n397;
wire            n398;
wire            n399;
wire            n400;
wire            n401;
wire            n402;
wire            n403;
wire            n404;
wire            n405;
wire            n406;
wire            n407;
wire            n408;
wire            n409;
wire            n410;
wire            n411;
wire            n412;
wire            n413;
wire            n414;
wire            n415;
wire            n416;
wire            n417;
wire            n418;
wire            n419;
wire            n420;
wire            n421;
wire            n422;
wire            n423;
wire            n424;
wire            n425;
wire            n426;
wire            n427;
wire            n428;
wire            n429;
wire            n430;
wire            n431;
wire            n432;
wire            n433;
wire            n434;
wire            n435;
wire            n436;
wire            n437;
wire            n438;
wire            n439;
wire            n440;
wire            n441;
wire            n442;
wire            n443;
wire            n444;
wire            n445;
wire            n446;
wire            n447;
wire            n448;
wire            n449;
wire            n450;
wire            n451;
wire            n452;
wire            n453;
wire            n454;
wire            n455;
wire            n456;
wire            n457;
wire            n458;
wire            n459;
wire            n460;
wire            n461;
wire            n462;
wire            n463;
wire            n464;
wire            n465;
wire            n466;
wire            n467;
wire            n468;
wire            n469;
wire            n470;
wire            n471;
wire            n472;
wire            n473;
wire            n474;
wire            n475;
wire            n476;
wire            n477;
wire            n478;
wire            n479;
wire            n480;
wire            n481;
wire            n482;
wire            n483;
wire            n484;
wire            n485;
wire            n486;
wire            n487;
wire            n488;
wire            n489;
wire            n490;
wire            n491;
wire            n492;
wire            n493;
wire            n494;
wire            n495;
wire            n496;
wire            n497;
wire            n498;
wire            n499;
wire            n500;
wire            n501;
wire            n502;
wire            n503;
wire            n504;
wire            n505;
wire            n506;
wire            n507;
wire            n508;
wire            n509;
wire            n510;
wire            n511;
wire            n512;
wire            n513;
wire            n514;
wire            n515;
wire            n516;
wire            n517;
wire            n518;
wire            n519;
wire            n520;
wire            n521;
wire            n522;
wire            n523;
wire            n524;
wire            n525;
wire            n526;
wire            n527;
wire            n528;
wire            n529;
wire            n530;
wire            n531;
wire            n532;
wire            n533;
wire            n534;
wire            n535;
wire            n536;
wire            n537;
wire            n538;
wire            n539;
wire            n540;
wire            n541;
wire            n542;
wire            n543;
wire            n544;
wire            n545;
wire            n546;
wire            n547;
wire            n548;
wire            n549;
wire            n550;
wire            n551;
wire            n552;
wire            n553;
wire            n554;
wire            n555;
wire            n556;
wire     [31:0] n557;
wire     [31:0] n558;
wire     [31:0] n559;
wire     [31:0] n560;
wire     [31:0] n561;
wire     [31:0] n562;
wire     [31:0] n563;
wire     [31:0] n564;
wire     [31:0] n565;
wire     [31:0] n566;
wire     [31:0] n567;
wire     [31:0] n568__choose_except;
wire     [31:0] n569;
wire     [31:0] n570;
wire            n571;
wire     [31:0] n572;
wire            n573;
wire            n574;
wire            n575;
wire            n576;
wire            n577;
wire            n578;
wire            n579;
wire            n580;
wire            n581;
wire            n582;
wire      [1:0] n583;
wire            n584;
wire      [1:0] n585;
wire            n586;
wire      [1:0] n587;
wire      [1:0] n588;
wire      [1:0] n589;
wire      [1:0] n590;
wire      [1:0] n591;
wire            n592;
wire            n593;
wire            n594;
wire            n595;
wire            n596;
wire            n597;
wire            n598;
wire            n599;
wire            n600;
wire            n601;
wire            n602;
wire            n603;
wire            n604;
wire            n605;
wire            n606;
wire            n607;
wire     [31:0] n608;
wire            n609;
wire            n610;
wire            n611;
wire            n612;
wire            n613;
wire            n614;
wire            n615;
wire            n616;
wire            n617;
wire            n618;
wire            n619;
wire            n620__take_int_or_expt;
wire            n621;
wire     [31:0] n622;
wire     [31:0] n623;
wire            n624;
wire            n625;
wire            n626;
wire            n627;
wire            n628;
wire            n629;
wire            n630;
wire            n631;
wire            n632;
wire            n633;
wire            n634;
wire            n635;
wire            n636;
wire            n637;
wire            n638;
wire            n639;
wire            n640;
wire            n641;
wire            n642;
wire     [31:0] n643;
wire     [31:0] n644;
wire     [31:0] n645;
wire     [31:0] n646;
wire     [31:0] n647;
wire     [31:0] n648;
wire     [31:0] n649;
wire     [31:0] n650;
wire     [31:0] n651;
wire     [31:0] n652;
wire     [31:0] n653;
wire     [31:0] n654;
wire     [31:0] n655;
wire     [31:0] n656;
wire     [31:0] n657;
wire     [31:0] n658;
wire     [31:0] n659;
wire     [31:0] n660;
wire     [31:0] n661;
wire     [31:0] n662;
wire     [31:0] n663;
wire     [31:0] n664;
wire     [31:0] n665;
wire     [31:0] n666;
wire     [31:0] n667__exception_code;
wire     [31:0] n668;
wire     [31:0] n669;
wire     [31:0] n670;
wire     [31:0] n671;
wire     [31:0] n672;
wire     [31:0] n673;
wire     [31:0] n674;
wire     [31:0] n675;
wire     [31:0] n676;
wire     [31:0] n677;
wire     [31:0] n678;
wire     [31:0] n679;
wire            n680;
wire            n681;
wire            n682;
wire      [1:0] n683;
wire      [1:0] n684;
wire            n685;
wire            n686;
wire            n687;
wire            n688;
wire            n689;
wire            n690;
wire            n691;
wire            n692;
wire            n693;
wire            n694;
wire            n695;
wire            n696;
wire            n697;
wire            n698;
wire            n699;
wire            n700;
wire            n701;
wire            n702;
wire            n703;
wire            n704;
wire            n705;
wire            n706;
wire            n707;
wire            n708;
wire            n709;
wire            n710;
wire            n711;
wire            n712;
wire            n713;
wire            n714;
wire            n715;
wire            n716;
wire            n717;
wire            n718;
wire            n719;
wire            n720;
wire      [1:0] n721;
wire      [2:0] n722;
wire      [3:0] n723;
wire      [4:0] n724;
wire      [5:0] n725;
wire      [6:0] n726;
wire      [7:0] n727;
wire      [8:0] n728;
wire     [10:0] n729;
wire     [12:0] n730;
wire     [31:0] n731;
wire     [31:0] n732;
wire     [31:0] n733;
wire     [31:0] n734;
wire     [31:0] n735;
wire     [31:0] n736;
wire     [31:0] n737;
wire     [31:0] n738;
wire     [31:0] n739;
wire      [6:0] n740;
wire            n741;
wire      [2:0] n742;
wire            n743;
wire            n744;
wire      [4:0] n745;
wire            n746;
wire            n747;
wire            n748;
wire            n749;
wire            n750;
wire            n751;
wire            n752;
wire            n753;
wire            n754;
wire            n755;
wire            n756;
wire            n757;
wire            n758;
wire            n759;
wire            n760;
wire            n761;
wire            n762;
wire            n763;
wire            n764;
wire            n765;
wire            n766;
wire            n767;
wire            n768;
wire            n769;
wire            n770;
wire            n771;
wire            n772;
wire            n773;
wire            n774;
wire            n775;
wire            n776;
wire     [31:0] n777;
wire     [31:0] n778;
wire     [31:0] n779;
wire     [31:0] n780;
wire     [31:0] n781;
wire     [31:0] n782;
wire     [31:0] n783;
wire     [31:0] n784;
wire     [31:0] n785;
wire     [31:0] n786;
wire     [31:0] n787;
wire     [31:0] n788;
wire     [31:0] n789;
wire     [31:0] n790;
wire     [31:0] n791;
wire     [31:0] n792;
wire     [31:0] n793;
wire     [31:0] n794;
wire     [31:0] n795;
wire     [31:0] n796;
wire     [31:0] n797;
wire     [31:0] n798;
wire     [31:0] n799;
wire     [31:0] n800;
wire     [31:0] n801;
wire     [31:0] n802;
wire     [31:0] n803;
wire     [31:0] n804;
wire     [31:0] n805;
wire     [31:0] n806;
wire     [31:0] n807;
wire     [11:0] n808;
wire     [31:0] n809;
wire     [31:0] n810;
wire     [31:0] n811;
wire            n812;
wire            n813;
wire      [7:0] n814;
wire            n815;
wire      [9:0] n816;
wire     [10:0] n817;
wire     [11:0] n818;
wire     [19:0] n819;
wire     [20:0] n820;
wire     [31:0] n821;
wire     [31:0] n822;
wire            n823;
wire            n824;
wire            n825;
wire      [4:0] n826;
wire            n827;
wire            n828;
wire            n829;
wire            n830;
wire            n831;
wire            n832;
wire            n833;
wire            n834;
wire            n835;
wire            n836;
wire            n837;
wire            n838;
wire            n839;
wire            n840;
wire            n841;
wire            n842;
wire            n843;
wire            n844;
wire            n845;
wire            n846;
wire            n847;
wire            n848;
wire            n849;
wire            n850;
wire            n851;
wire            n852;
wire            n853;
wire            n854;
wire            n855;
wire            n856;
wire            n857;
wire     [31:0] n858;
wire     [31:0] n859;
wire     [31:0] n860;
wire     [31:0] n861;
wire     [31:0] n862;
wire     [31:0] n863;
wire     [31:0] n864;
wire     [31:0] n865;
wire     [31:0] n866;
wire     [31:0] n867;
wire     [31:0] n868;
wire     [31:0] n869;
wire     [31:0] n870;
wire     [31:0] n871;
wire     [31:0] n872;
wire     [31:0] n873;
wire     [31:0] n874;
wire     [31:0] n875;
wire     [31:0] n876;
wire     [31:0] n877;
wire     [31:0] n878;
wire     [31:0] n879;
wire     [31:0] n880;
wire     [31:0] n881;
wire     [31:0] n882;
wire     [31:0] n883;
wire     [31:0] n884;
wire     [31:0] n885;
wire     [31:0] n886;
wire     [31:0] n887;
wire     [31:0] n888;
wire            n889;
wire            n890;
wire      [5:0] n891;
wire      [3:0] n892;
wire      [4:0] n893;
wire     [10:0] n894;
wire     [11:0] n895;
wire     [12:0] n896;
wire     [31:0] n897;
wire     [31:0] n898;
wire     [31:0] n899;
wire     [31:0] n900;
wire            n901;
wire            n902;
wire            n903;
wire     [31:0] n904;
wire            n905;
wire            n906;
wire            n907;
wire     [31:0] n908;
wire            n909;
wire            n910;
wire            n911;
wire     [31:0] n912;
wire            n913;
wire            n914;
wire            n915;
wire     [31:0] n916;
wire            n917;
wire            n918;
wire     [31:0] n919;
wire            n920;
wire            n921;
wire      [6:0] n922;
wire            n923;
wire            n924;
wire            n925;
wire            n926;
wire            n927;
wire            n928;
wire            n929;
wire            n930;
wire            n931;
wire            n932;
wire            n933;
wire            n934;
wire            n935;
wire            n936;
wire            n937;
wire            n938;
wire            n939;
wire            n940;
wire            n941;
wire            n942;
wire            n943;
wire            n944;
wire            n945;
wire            n946;
wire            n947;
wire            n948;
wire            n949;
wire            n950;
wire            n951;
wire            n952;
wire            n953;
wire            n954;
wire            n955;
wire            n956;
wire            n957;
wire            n958;
wire            n959;
wire            n960;
wire            n961;
wire            n962;
wire            n963;
wire            n964;
wire            n965;
wire            n966;
wire            n967;
wire            n968;
wire            n969;
wire            n970;
wire            n971;
wire            n972;
wire            n973;
wire            n974;
wire            n975;
wire            n976;
wire            n977;
wire            n978;
wire            n979;
wire            n980;
wire            n981;
wire            n982;
wire            n983;
wire            n984;
wire            n985;
wire            n986;
wire            n987;
wire            n988;
wire            n989;
wire            n990;
wire            n991;
wire            n992;
wire            n993;
wire            n994;
wire            n995;
wire     [31:0] n996;
wire     [31:0] n997;
wire     [31:0] n998;
wire     [31:0] n999;
wire     [31:0] n1000;
wire     [31:0] n1001;
wire     [31:0] n1002;
wire     [31:0] n1003;
wire     [31:0] n1004;
wire     [31:0] n1005;
wire     [31:0] n1006;
wire     [31:0] n1007;
wire            n1008;
wire     [31:0] n1009;
wire     [31:0] n1010;
wire            n1011;
wire     [31:0] n1012;
wire     [31:0] n1013;
wire     [31:0] n1014;
wire     [31:0] n1015;
wire     [31:0] n1016;
wire     [31:0] n1017;
wire     [31:0] n1018;
wire     [31:0] n1019;
wire     [31:0] n1020;
wire      [4:0] n1021;
wire            n1022;
wire      [4:0] n1023;
wire     [31:0] n1024;
wire     [31:0] n1025;
wire     [31:0] n1026;
wire     [31:0] n1027;
wire     [31:0] n1028;
wire     [31:0] n1029;
wire     [31:0] n1030;
wire     [31:0] n1031;
wire     [31:0] n1032;
wire     [31:0] n1033;
wire     [31:0] n1034;
wire     [31:0] n1035;
wire     [31:0] n1036;
wire     [31:0] n1037;
wire     [31:0] n1038;
wire     [31:0] n1039;
wire     [31:0] n1040;
wire     [31:0] n1041;
wire     [31:0] n1042;
wire     [31:0] n1043;
wire     [31:0] n1044;
wire     [31:0] n1045;
wire     [31:0] n1046;
wire     [31:0] n1047;
wire     [31:0] n1048;
wire     [31:0] n1049;
wire     [31:0] n1050;
wire     [31:0] n1051;
wire     [31:0] n1052;
wire     [31:0] n1053;
wire     [31:0] n1054;
wire     [31:0] n1055;
wire     [31:0] n1056;
wire     [31:0] n1057;
wire     [31:0] n1058;
wire     [31:0] n1059;
wire            n1060;
wire     [31:0] n1061;
wire     [31:0] n1062;
wire            n1063;
wire     [31:0] n1064;
wire     [31:0] n1065;
wire     [31:0] n1066;
wire     [31:0] n1067;
wire            n1068;
wire     [31:0] n1069;
wire     [19:0] n1070;
wire     [31:0] n1071;
wire     [31:0] n1072;
wire     [31:0] n1073;
wire     [31:0] n1074;
wire      [1:0] n1075;
wire            n1076;
wire     [29:0] n1077;
wire     [31:0] n1078;
wire     [31:0] n1081;
wire     [15:0] n1082;
wire     [31:0] n1083;
wire            n1084;
wire      [7:0] n1085;
wire     [31:0] n1086;
wire            n1087;
wire     [15:0] n1088;
wire     [31:0] n1089;
wire            n1090;
wire      [7:0] n1091;
wire     [31:0] n1092;
wire     [31:0] n1093;
wire     [31:0] n1094;
wire     [31:0] n1095;
wire     [31:0] n1096;
wire     [31:0] n1097;
wire     [31:0] n1098;
wire      [7:0] n1099;
wire     [31:0] n1100;
wire      [7:0] n1101;
wire     [31:0] n1102;
wire     [31:0] n1103;
wire     [31:0] n1104;
wire     [31:0] n1105;
wire     [31:0] n1106;
wire     [31:0] n1107;
wire     [31:0] n1108;
wire     [31:0] n1109;
wire     [31:0] n1110;
wire     [31:0] n1111;
wire     [31:0] n1112;
wire     [31:0] n1113;
wire     [31:0] n1114;
wire     [31:0] n1115;
wire     [31:0] n1116;
wire     [31:0] n1117;
wire     [31:0] n1118;
wire     [31:0] n1119;
wire     [31:0] n1120;
wire     [31:0] n1121;
wire     [31:0] n1122;
wire     [31:0] n1123;
wire     [31:0] n1124;
wire     [31:0] n1125;
wire     [31:0] n1126;
wire     [31:0] n1127;
wire     [31:0] n1128;
wire     [31:0] n1129;
wire     [31:0] n1130;
wire     [31:0] n1131;
wire     [31:0] n1132;
wire     [31:0] n1133;
wire     [31:0] n1134;
wire     [31:0] n1135;
wire     [31:0] n1136;
wire     [31:0] n1137;
wire     [31:0] n1138;
wire     [31:0] n1139;
wire     [31:0] n1140;
wire     [31:0] n1141;
wire     [31:0] n1142;
wire     [31:0] n1143;
wire     [31:0] n1144;
wire     [31:0] n1145;
wire     [31:0] n1146;
wire     [31:0] n1147;
wire     [31:0] n1148;
wire     [31:0] n1149;
wire     [31:0] n1150;
wire     [31:0] n1151;
wire            n1152;
wire     [31:0] n1153;
wire     [31:0] n1154;
wire     [31:0] n1155;
wire     [31:0] n1156;
wire     [31:0] n1157;
wire     [31:0] n1158;
wire     [31:0] n1159;
wire     [31:0] n1160;
wire     [31:0] n1161;
wire     [31:0] n1162;
wire     [31:0] n1163;
wire     [31:0] n1164;
wire     [31:0] n1165;
wire     [31:0] n1166;
wire     [31:0] n1167;
wire     [31:0] n1168;
wire     [31:0] n1169;
wire     [31:0] n1170;
wire     [31:0] n1171;
wire     [31:0] n1172;
wire     [31:0] n1173;
wire     [31:0] n1174;
wire     [31:0] n1175;
wire     [31:0] n1176;
wire     [31:0] n1177;
wire     [31:0] n1178;
wire     [31:0] n1179;
wire     [31:0] n1180;
wire     [31:0] n1181;
wire     [31:0] n1182;
wire     [31:0] n1183;
wire     [31:0] n1184;
wire     [31:0] n1185;
wire     [31:0] n1186;
wire     [31:0] n1187;
wire     [31:0] n1188;
wire     [31:0] n1189;
wire     [31:0] n1190;
wire     [31:0] n1191;
wire     [31:0] n1192;
wire     [31:0] n1193;
wire     [31:0] n1194;
wire     [31:0] n1195;
wire     [31:0] n1196;
wire     [31:0] n1197;
wire     [31:0] n1198;
wire     [31:0] n1199;
wire     [31:0] n1200;
wire     [31:0] n1201;
wire     [31:0] n1202;
wire     [31:0] n1203;
wire     [31:0] n1204;
wire     [31:0] n1205;
wire     [31:0] n1206;
wire     [31:0] n1207;
wire     [31:0] n1208;
wire            n1209;
wire     [31:0] n1210;
wire     [31:0] n1211;
wire     [31:0] n1212;
wire     [31:0] n1213;
wire     [31:0] n1214;
wire     [31:0] n1215;
wire     [31:0] n1216;
wire     [31:0] n1217;
wire     [31:0] n1218;
wire     [31:0] n1219;
wire     [31:0] n1220;
wire     [31:0] n1221;
wire     [31:0] n1222;
wire     [31:0] n1223;
wire     [31:0] n1224;
wire     [31:0] n1225;
wire     [31:0] n1226;
wire     [31:0] n1227;
wire     [31:0] n1228;
wire     [31:0] n1229;
wire     [31:0] n1230;
wire     [31:0] n1231;
wire     [31:0] n1232;
wire     [31:0] n1233;
wire     [31:0] n1234;
wire     [31:0] n1235;
wire     [31:0] n1236;
wire     [31:0] n1237;
wire     [31:0] n1238;
wire     [31:0] n1239;
wire     [31:0] n1240;
wire     [31:0] n1241;
wire     [31:0] n1242;
wire     [31:0] n1243;
wire     [31:0] n1244;
wire     [31:0] n1245;
wire     [31:0] n1246;
wire     [31:0] n1247;
wire     [31:0] n1248;
wire     [31:0] n1249;
wire     [31:0] n1250;
wire     [31:0] n1251;
wire     [31:0] n1252;
wire     [31:0] n1253;
wire     [31:0] n1254;
wire     [31:0] n1255;
wire     [31:0] n1256;
wire     [31:0] n1257;
wire     [31:0] n1258;
wire     [31:0] n1259;
wire     [31:0] n1260;
wire     [31:0] n1261;
wire     [31:0] n1262;
wire     [31:0] n1263;
wire     [31:0] n1264;
wire            n1265;
wire     [31:0] n1266;
wire     [31:0] n1267;
wire     [31:0] n1268;
wire     [31:0] n1269;
wire     [31:0] n1270;
wire     [31:0] n1271;
wire     [31:0] n1272;
wire     [31:0] n1273;
wire     [31:0] n1274;
wire     [31:0] n1275;
wire     [31:0] n1276;
wire     [31:0] n1277;
wire     [31:0] n1278;
wire     [31:0] n1279;
wire     [31:0] n1280;
wire     [31:0] n1281;
wire            n1282;
wire     [31:0] n1283;
wire     [31:0] n1284;
wire     [31:0] n1285;
wire     [31:0] n1286;
wire     [31:0] n1287;
wire     [31:0] n1288;
wire     [31:0] n1289;
wire     [31:0] n1290;
wire     [31:0] n1291;
wire     [31:0] n1292;
wire     [31:0] n1293;
wire     [31:0] n1294;
wire     [31:0] n1295;
wire     [31:0] n1296;
wire     [31:0] n1297;
wire     [31:0] n1298;
wire     [31:0] n1299;
wire     [31:0] n1300;
wire     [31:0] n1301;
wire     [31:0] n1302;
wire     [31:0] n1303;
wire     [31:0] n1304;
wire     [31:0] n1305;
wire     [31:0] n1306;
wire     [31:0] n1307;
wire     [31:0] n1308;
wire     [31:0] n1309;
wire     [31:0] n1310;
wire     [31:0] n1311;
wire     [31:0] n1312;
wire     [31:0] n1313;
wire     [31:0] n1314;
wire     [31:0] n1315;
wire     [31:0] n1316;
wire     [31:0] n1317;
wire     [31:0] n1318;
wire     [31:0] n1319;
wire     [31:0] n1320;
wire     [31:0] n1321;
wire     [31:0] n1322;
wire            n1323;
wire     [31:0] n1324;
wire     [31:0] n1325;
wire     [31:0] n1326;
wire     [31:0] n1327;
wire     [31:0] n1328;
wire     [31:0] n1329;
wire     [31:0] n1330;
wire     [31:0] n1331;
wire     [31:0] n1332;
wire     [31:0] n1333;
wire     [31:0] n1334;
wire     [31:0] n1335;
wire     [31:0] n1336;
wire     [31:0] n1337;
wire     [31:0] n1338;
wire     [31:0] n1339;
wire     [31:0] n1340;
wire     [31:0] n1341;
wire            n1342;
wire     [31:0] n1343;
wire     [31:0] n1344;
wire     [31:0] n1345;
wire     [31:0] n1346;
wire     [31:0] n1347;
wire     [31:0] n1348;
wire     [31:0] n1349;
wire     [31:0] n1350;
wire     [31:0] n1351;
wire     [31:0] n1352;
wire     [31:0] n1353;
wire     [31:0] n1354;
wire     [31:0] n1355;
wire     [31:0] n1356;
wire     [31:0] n1357;
wire     [31:0] n1358;
wire     [31:0] n1359;
wire     [31:0] n1360;
wire     [31:0] n1361;
wire     [31:0] n1362;
wire     [31:0] n1363;
wire     [31:0] n1364;
wire     [31:0] n1365;
wire     [31:0] n1366;
wire     [31:0] n1367;
wire     [31:0] n1368;
wire     [31:0] n1369;
wire     [31:0] n1370;
wire     [31:0] n1371;
wire     [31:0] n1372;
wire     [31:0] n1373;
wire     [31:0] n1374;
wire     [31:0] n1375;
wire     [31:0] n1376;
wire     [31:0] n1377;
wire     [31:0] n1378;
wire     [31:0] n1379;
wire     [31:0] n1380;
wire     [31:0] n1381;
wire            n1382;
wire     [31:0] n1383;
wire     [31:0] n1384;
wire     [31:0] n1385;
wire     [31:0] n1386;
wire     [31:0] n1387;
wire     [31:0] n1388;
wire     [31:0] n1389;
wire     [31:0] n1390;
wire     [31:0] n1391;
wire     [31:0] n1392;
wire     [31:0] n1393;
wire     [31:0] n1394;
wire     [31:0] n1395;
wire     [31:0] n1396;
wire     [31:0] n1397;
wire     [31:0] n1398;
wire     [31:0] n1399;
wire     [31:0] n1400;
wire     [31:0] n1401;
wire     [31:0] n1402;
wire     [31:0] n1403;
wire     [31:0] n1404;
wire     [31:0] n1405;
wire     [31:0] n1406;
wire     [31:0] n1407;
wire     [31:0] n1408;
wire     [31:0] n1409;
wire     [31:0] n1410;
wire     [31:0] n1411;
wire     [31:0] n1412;
wire     [31:0] n1413;
wire     [31:0] n1414;
wire     [31:0] n1415;
wire     [31:0] n1416;
wire     [31:0] n1417;
wire     [31:0] n1418;
wire     [31:0] n1419;
wire     [31:0] n1420;
wire     [31:0] n1421;
wire     [31:0] n1422;
wire     [31:0] n1423;
wire     [31:0] n1424;
wire     [31:0] n1425;
wire     [31:0] n1426;
wire     [31:0] n1427;
wire     [31:0] n1428;
wire     [31:0] n1429;
wire     [31:0] n1430;
wire     [31:0] n1431;
wire     [31:0] n1432;
wire     [31:0] n1433;
wire     [31:0] n1434;
wire     [31:0] n1435;
wire     [31:0] n1436;
wire     [31:0] n1437;
wire            n1438;
wire     [31:0] n1439;
wire     [31:0] n1440;
wire     [31:0] n1441;
wire     [31:0] n1442;
wire     [31:0] n1443;
wire     [31:0] n1444;
wire     [31:0] n1445;
wire     [31:0] n1446;
wire     [31:0] n1447;
wire     [31:0] n1448;
wire     [31:0] n1449;
wire     [31:0] n1450;
wire     [31:0] n1451;
wire     [31:0] n1452;
wire     [31:0] n1453;
wire     [31:0] n1454;
wire     [31:0] n1455;
wire     [31:0] n1456;
wire     [31:0] n1457;
wire     [31:0] n1458;
wire     [31:0] n1459;
wire     [31:0] n1460;
wire     [31:0] n1461;
wire     [31:0] n1462;
wire     [31:0] n1463;
wire     [31:0] n1464;
wire     [31:0] n1465;
wire     [31:0] n1466;
wire     [31:0] n1467;
wire     [31:0] n1468;
wire     [31:0] n1469;
wire     [31:0] n1470;
wire     [31:0] n1471;
wire     [31:0] n1472;
wire     [31:0] n1473;
wire     [31:0] n1474;
wire     [31:0] n1475;
wire     [31:0] n1476;
wire     [31:0] n1477;
wire     [31:0] n1478;
wire     [31:0] n1479;
wire     [31:0] n1480;
wire     [31:0] n1481;
wire     [31:0] n1482;
wire     [31:0] n1483;
wire     [31:0] n1484;
wire     [31:0] n1485;
wire     [31:0] n1486;
wire     [31:0] n1487;
wire     [31:0] n1488;
wire     [31:0] n1489;
wire     [31:0] n1490;
wire     [31:0] n1491;
wire     [31:0] n1492;
wire     [31:0] n1493;
wire     [31:0] n1494;
wire            n1495;
wire     [31:0] n1496;
wire     [31:0] n1497;
wire     [31:0] n1498;
wire     [31:0] n1499;
wire     [31:0] n1500;
wire     [31:0] n1501;
wire     [31:0] n1502;
wire     [31:0] n1503;
wire     [31:0] n1504;
wire     [31:0] n1505;
wire     [31:0] n1506;
wire     [31:0] n1507;
wire     [31:0] n1508;
wire     [31:0] n1509;
wire     [31:0] n1510;
wire     [31:0] n1511;
wire     [31:0] n1512;
wire     [31:0] n1513;
wire     [31:0] n1514;
wire     [31:0] n1515;
wire     [31:0] n1516;
wire     [31:0] n1517;
wire     [31:0] n1518;
wire     [31:0] n1519;
wire     [31:0] n1520;
wire     [31:0] n1521;
wire     [31:0] n1522;
wire     [31:0] n1523;
wire     [31:0] n1524;
wire     [31:0] n1525;
wire     [31:0] n1526;
wire     [31:0] n1527;
wire     [31:0] n1528;
wire     [31:0] n1529;
wire     [31:0] n1530;
wire     [31:0] n1531;
wire     [31:0] n1532;
wire     [31:0] n1533;
wire     [31:0] n1534;
wire     [31:0] n1535;
wire     [31:0] n1536;
wire     [31:0] n1537;
wire     [31:0] n1538;
wire     [31:0] n1539;
wire     [31:0] n1540;
wire     [31:0] n1541;
wire     [31:0] n1542;
wire     [31:0] n1543;
wire     [31:0] n1544;
wire     [31:0] n1545;
wire     [31:0] n1546;
wire     [31:0] n1547;
wire     [31:0] n1548;
wire     [31:0] n1549;
wire     [31:0] n1550;
wire            n1551;
wire     [31:0] n1552;
wire     [31:0] n1553;
wire     [31:0] n1554;
wire     [31:0] n1555;
wire     [31:0] n1556;
wire     [31:0] n1557;
wire     [31:0] n1558;
wire     [31:0] n1559;
wire     [31:0] n1560;
wire     [31:0] n1561;
wire     [31:0] n1562;
wire     [31:0] n1563;
wire     [31:0] n1564;
wire     [31:0] n1565;
wire     [31:0] n1566;
wire     [31:0] n1567;
wire     [31:0] n1568;
wire     [31:0] n1569;
wire     [31:0] n1570;
wire     [31:0] n1571;
wire     [31:0] n1572;
wire     [31:0] n1573;
wire     [31:0] n1574;
wire     [31:0] n1575;
wire     [31:0] n1576;
wire     [31:0] n1577;
wire     [31:0] n1578;
wire     [31:0] n1579;
wire     [31:0] n1580;
wire     [31:0] n1581;
wire     [31:0] n1582;
wire     [31:0] n1583;
wire     [31:0] n1584;
wire     [31:0] n1585;
wire     [31:0] n1586;
wire     [31:0] n1587;
wire     [31:0] n1588;
wire     [31:0] n1589;
wire     [31:0] n1590;
wire     [31:0] n1591;
wire     [31:0] n1592;
wire     [31:0] n1593;
wire     [31:0] n1594;
wire     [31:0] n1595;
wire     [31:0] n1596;
wire     [31:0] n1597;
wire     [31:0] n1598;
wire     [31:0] n1599;
wire     [31:0] n1600;
wire     [31:0] n1601;
wire     [31:0] n1602;
wire     [31:0] n1603;
wire     [31:0] n1604;
wire     [31:0] n1605;
wire     [31:0] n1606;
wire            n1607;
wire     [31:0] n1608;
wire     [31:0] n1609;
wire     [31:0] n1610;
wire     [31:0] n1611;
wire     [31:0] n1612;
wire     [31:0] n1613;
wire     [31:0] n1614;
wire     [31:0] n1615;
wire     [31:0] n1616;
wire     [31:0] n1617;
wire     [31:0] n1618;
wire     [31:0] n1619;
wire     [31:0] n1620;
wire     [31:0] n1621;
wire     [31:0] n1622;
wire     [31:0] n1623;
wire     [31:0] n1624;
wire     [31:0] n1625;
wire     [31:0] n1626;
wire     [31:0] n1627;
wire     [31:0] n1628;
wire     [31:0] n1629;
wire     [31:0] n1630;
wire     [31:0] n1631;
wire     [31:0] n1632;
wire     [31:0] n1633;
wire     [31:0] n1634;
wire     [31:0] n1635;
wire     [31:0] n1636;
wire     [31:0] n1637;
wire     [31:0] n1638;
wire     [31:0] n1639;
wire     [31:0] n1640;
wire     [31:0] n1641;
wire     [31:0] n1642;
wire     [31:0] n1643;
wire     [31:0] n1644;
wire     [31:0] n1645;
wire     [31:0] n1646;
wire     [31:0] n1647;
wire     [31:0] n1648;
wire     [31:0] n1649;
wire     [31:0] n1650;
wire     [31:0] n1651;
wire     [31:0] n1652;
wire     [31:0] n1653;
wire     [31:0] n1654;
wire     [31:0] n1655;
wire     [31:0] n1656;
wire     [31:0] n1657;
wire     [31:0] n1658;
wire     [31:0] n1659;
wire     [31:0] n1660;
wire     [31:0] n1661;
wire     [31:0] n1662;
wire            n1663;
wire     [31:0] n1664;
wire     [31:0] n1665;
wire     [31:0] n1666;
wire     [31:0] n1667;
wire     [31:0] n1668;
wire     [31:0] n1669;
wire     [31:0] n1670;
wire     [31:0] n1671;
wire     [31:0] n1672;
wire     [31:0] n1673;
wire     [31:0] n1674;
wire     [31:0] n1675;
wire     [31:0] n1676;
wire     [31:0] n1677;
wire     [31:0] n1678;
wire     [31:0] n1679;
wire     [31:0] n1680;
wire     [31:0] n1681;
wire     [31:0] n1682;
wire     [31:0] n1683;
wire     [31:0] n1684;
wire     [31:0] n1685;
wire     [31:0] n1686;
wire     [31:0] n1687;
wire     [31:0] n1688;
wire     [31:0] n1689;
wire     [31:0] n1690;
wire     [31:0] n1691;
wire     [31:0] n1692;
wire     [31:0] n1693;
wire     [31:0] n1694;
wire     [31:0] n1695;
wire     [31:0] n1696;
wire     [31:0] n1697;
wire     [31:0] n1698;
wire     [31:0] n1699;
wire     [31:0] n1700;
wire     [31:0] n1701;
wire     [31:0] n1702;
wire     [31:0] n1703;
wire     [31:0] n1704;
wire     [31:0] n1705;
wire     [31:0] n1706;
wire     [31:0] n1707;
wire     [31:0] n1708;
wire     [31:0] n1709;
wire     [31:0] n1710;
wire     [31:0] n1711;
wire     [31:0] n1712;
wire     [31:0] n1713;
wire     [31:0] n1714;
wire     [31:0] n1715;
wire     [31:0] n1716;
wire     [31:0] n1717;
wire     [31:0] n1718;
wire            n1719;
wire     [31:0] n1720;
wire     [31:0] n1721;
wire     [31:0] n1722;
wire     [31:0] n1723;
wire     [31:0] n1724;
wire     [31:0] n1725;
wire     [31:0] n1726;
wire     [31:0] n1727;
wire     [31:0] n1728;
wire     [31:0] n1729;
wire     [31:0] n1730;
wire     [31:0] n1731;
wire     [31:0] n1732;
wire     [31:0] n1733;
wire     [31:0] n1734;
wire     [31:0] n1735;
wire     [31:0] n1736;
wire     [31:0] n1737;
wire     [31:0] n1738;
wire     [31:0] n1739;
wire     [31:0] n1740;
wire     [31:0] n1741;
wire     [31:0] n1742;
wire     [31:0] n1743;
wire     [31:0] n1744;
wire     [31:0] n1745;
wire     [31:0] n1746;
wire     [31:0] n1747;
wire     [31:0] n1748;
wire     [31:0] n1749;
wire     [31:0] n1750;
wire     [31:0] n1751;
wire     [31:0] n1752;
wire     [31:0] n1753;
wire     [31:0] n1754;
wire     [31:0] n1755;
wire     [31:0] n1756;
wire     [31:0] n1757;
wire     [31:0] n1758;
wire     [31:0] n1759;
wire     [31:0] n1760;
wire     [31:0] n1761;
wire     [31:0] n1762;
wire     [31:0] n1763;
wire     [31:0] n1764;
wire     [31:0] n1765;
wire     [31:0] n1766;
wire     [31:0] n1767;
wire     [31:0] n1768;
wire     [31:0] n1769;
wire     [31:0] n1770;
wire     [31:0] n1771;
wire     [31:0] n1772;
wire     [31:0] n1773;
wire     [31:0] n1774;
wire            n1775;
wire     [31:0] n1776;
wire     [31:0] n1777;
wire     [31:0] n1778;
wire     [31:0] n1779;
wire     [31:0] n1780;
wire     [31:0] n1781;
wire     [31:0] n1782;
wire     [31:0] n1783;
wire     [31:0] n1784;
wire     [31:0] n1785;
wire     [31:0] n1786;
wire     [31:0] n1787;
wire     [31:0] n1788;
wire     [31:0] n1789;
wire     [31:0] n1790;
wire     [31:0] n1791;
wire     [31:0] n1792;
wire     [31:0] n1793;
wire     [31:0] n1794;
wire     [31:0] n1795;
wire     [31:0] n1796;
wire     [31:0] n1797;
wire     [31:0] n1798;
wire     [31:0] n1799;
wire     [31:0] n1800;
wire     [31:0] n1801;
wire     [31:0] n1802;
wire     [31:0] n1803;
wire     [31:0] n1804;
wire     [31:0] n1805;
wire     [31:0] n1806;
wire     [31:0] n1807;
wire     [31:0] n1808;
wire     [31:0] n1809;
wire     [31:0] n1810;
wire     [31:0] n1811;
wire     [31:0] n1812;
wire     [31:0] n1813;
wire     [31:0] n1814;
wire     [31:0] n1815;
wire     [31:0] n1816;
wire     [31:0] n1817;
wire     [31:0] n1818;
wire     [31:0] n1819;
wire     [31:0] n1820;
wire     [31:0] n1821;
wire     [31:0] n1822;
wire     [31:0] n1823;
wire     [31:0] n1824;
wire     [31:0] n1825;
wire     [31:0] n1826;
wire     [31:0] n1827;
wire     [31:0] n1828;
wire     [31:0] n1829;
wire     [31:0] n1830;
wire            n1831;
wire     [31:0] n1832;
wire     [31:0] n1833;
wire     [31:0] n1834;
wire     [31:0] n1835;
wire     [31:0] n1836;
wire     [31:0] n1837;
wire     [31:0] n1838;
wire     [31:0] n1839;
wire     [31:0] n1840;
wire     [31:0] n1841;
wire     [31:0] n1842;
wire     [31:0] n1843;
wire     [31:0] n1844;
wire     [31:0] n1845;
wire     [31:0] n1846;
wire     [31:0] n1847;
wire     [31:0] n1848;
wire     [31:0] n1849;
wire     [31:0] n1850;
wire     [31:0] n1851;
wire     [31:0] n1852;
wire     [31:0] n1853;
wire     [31:0] n1854;
wire     [31:0] n1855;
wire     [31:0] n1856;
wire     [31:0] n1857;
wire     [31:0] n1858;
wire     [31:0] n1859;
wire     [31:0] n1860;
wire     [31:0] n1861;
wire     [31:0] n1862;
wire     [31:0] n1863;
wire     [31:0] n1864;
wire     [31:0] n1865;
wire     [31:0] n1866;
wire     [31:0] n1867;
wire     [31:0] n1868;
wire     [31:0] n1869;
wire     [31:0] n1870;
wire     [31:0] n1871;
wire     [31:0] n1872;
wire     [31:0] n1873;
wire     [31:0] n1874;
wire     [31:0] n1875;
wire     [31:0] n1876;
wire     [31:0] n1877;
wire     [31:0] n1878;
wire     [31:0] n1879;
wire     [31:0] n1880;
wire     [31:0] n1881;
wire     [31:0] n1882;
wire     [31:0] n1883;
wire     [31:0] n1884;
wire     [31:0] n1885;
wire     [31:0] n1886;
wire            n1887;
wire     [31:0] n1888;
wire     [31:0] n1889;
wire     [31:0] n1890;
wire     [31:0] n1891;
wire     [31:0] n1892;
wire     [31:0] n1893;
wire     [31:0] n1894;
wire     [31:0] n1895;
wire     [31:0] n1896;
wire     [31:0] n1897;
wire     [31:0] n1898;
wire     [31:0] n1899;
wire     [31:0] n1900;
wire     [31:0] n1901;
wire     [31:0] n1902;
wire     [31:0] n1903;
wire     [31:0] n1904;
wire     [31:0] n1905;
wire     [31:0] n1906;
wire     [31:0] n1907;
wire     [31:0] n1908;
wire     [31:0] n1909;
wire     [31:0] n1910;
wire     [31:0] n1911;
wire     [31:0] n1912;
wire     [31:0] n1913;
wire     [31:0] n1914;
wire     [31:0] n1915;
wire     [31:0] n1916;
wire     [31:0] n1917;
wire     [31:0] n1918;
wire     [31:0] n1919;
wire     [31:0] n1920;
wire     [31:0] n1921;
wire     [31:0] n1922;
wire     [31:0] n1923;
wire     [31:0] n1924;
wire     [31:0] n1925;
wire     [31:0] n1926;
wire     [31:0] n1927;
wire     [31:0] n1928;
wire     [31:0] n1929;
wire     [31:0] n1930;
wire     [31:0] n1931;
wire     [31:0] n1932;
wire     [31:0] n1933;
wire     [31:0] n1934;
wire     [31:0] n1935;
wire     [31:0] n1936;
wire     [31:0] n1937;
wire     [31:0] n1938;
wire     [31:0] n1939;
wire     [31:0] n1940;
wire     [31:0] n1941;
wire     [31:0] n1942;
wire            n1943;
wire     [31:0] n1944;
wire     [31:0] n1945;
wire     [31:0] n1946;
wire     [31:0] n1947;
wire     [31:0] n1948;
wire     [31:0] n1949;
wire     [31:0] n1950;
wire     [31:0] n1951;
wire     [31:0] n1952;
wire     [31:0] n1953;
wire     [31:0] n1954;
wire     [31:0] n1955;
wire     [31:0] n1956;
wire     [31:0] n1957;
wire     [31:0] n1958;
wire     [31:0] n1959;
wire     [31:0] n1960;
wire     [31:0] n1961;
wire     [31:0] n1962;
wire     [31:0] n1963;
wire     [31:0] n1964;
wire     [31:0] n1965;
wire     [31:0] n1966;
wire     [31:0] n1967;
wire     [31:0] n1968;
wire     [31:0] n1969;
wire     [31:0] n1970;
wire     [31:0] n1971;
wire     [31:0] n1972;
wire     [31:0] n1973;
wire     [31:0] n1974;
wire     [31:0] n1975;
wire     [31:0] n1976;
wire     [31:0] n1977;
wire     [31:0] n1978;
wire     [31:0] n1979;
wire     [31:0] n1980;
wire     [31:0] n1981;
wire     [31:0] n1982;
wire     [31:0] n1983;
wire     [31:0] n1984;
wire     [31:0] n1985;
wire     [31:0] n1986;
wire     [31:0] n1987;
wire     [31:0] n1988;
wire     [31:0] n1989;
wire     [31:0] n1990;
wire     [31:0] n1991;
wire     [31:0] n1992;
wire     [31:0] n1993;
wire     [31:0] n1994;
wire     [31:0] n1995;
wire     [31:0] n1996;
wire     [31:0] n1997;
wire     [31:0] n1998;
wire            n1999;
wire     [31:0] n2000;
wire     [31:0] n2001;
wire     [31:0] n2002;
wire     [31:0] n2003;
wire     [31:0] n2004;
wire     [31:0] n2005;
wire     [31:0] n2006;
wire     [31:0] n2007;
wire     [31:0] n2008;
wire     [31:0] n2009;
wire     [31:0] n2010;
wire     [31:0] n2011;
wire     [31:0] n2012;
wire     [31:0] n2013;
wire     [31:0] n2014;
wire     [31:0] n2015;
wire     [31:0] n2016;
wire     [31:0] n2017;
wire     [31:0] n2018;
wire     [31:0] n2019;
wire     [31:0] n2020;
wire     [31:0] n2021;
wire     [31:0] n2022;
wire     [31:0] n2023;
wire     [31:0] n2024;
wire     [31:0] n2025;
wire     [31:0] n2026;
wire     [31:0] n2027;
wire     [31:0] n2028;
wire     [31:0] n2029;
wire     [31:0] n2030;
wire     [31:0] n2031;
wire     [31:0] n2032;
wire     [31:0] n2033;
wire     [31:0] n2034;
wire     [31:0] n2035;
wire     [31:0] n2036;
wire     [31:0] n2037;
wire     [31:0] n2038;
wire     [31:0] n2039;
wire     [31:0] n2040;
wire     [31:0] n2041;
wire     [31:0] n2042;
wire     [31:0] n2043;
wire     [31:0] n2044;
wire     [31:0] n2045;
wire     [31:0] n2046;
wire     [31:0] n2047;
wire     [31:0] n2048;
wire     [31:0] n2049;
wire     [31:0] n2050;
wire     [31:0] n2051;
wire     [31:0] n2052;
wire     [31:0] n2053;
wire     [31:0] n2054;
wire            n2055;
wire     [31:0] n2056;
wire     [31:0] n2057;
wire     [31:0] n2058;
wire     [31:0] n2059;
wire     [31:0] n2060;
wire     [31:0] n2061;
wire     [31:0] n2062;
wire     [31:0] n2063;
wire     [31:0] n2064;
wire     [31:0] n2065;
wire     [31:0] n2066;
wire     [31:0] n2067;
wire     [31:0] n2068;
wire     [31:0] n2069;
wire     [31:0] n2070;
wire     [31:0] n2071;
wire     [31:0] n2072;
wire     [31:0] n2073;
wire     [31:0] n2074;
wire     [31:0] n2075;
wire     [31:0] n2076;
wire     [31:0] n2077;
wire     [31:0] n2078;
wire     [31:0] n2079;
wire     [31:0] n2080;
wire     [31:0] n2081;
wire     [31:0] n2082;
wire     [31:0] n2083;
wire     [31:0] n2084;
wire     [31:0] n2085;
wire     [31:0] n2086;
wire     [31:0] n2087;
wire     [31:0] n2088;
wire     [31:0] n2089;
wire     [31:0] n2090;
wire     [31:0] n2091;
wire     [31:0] n2092;
wire     [31:0] n2093;
wire     [31:0] n2094;
wire     [31:0] n2095;
wire     [31:0] n2096;
wire     [31:0] n2097;
wire     [31:0] n2098;
wire     [31:0] n2099;
wire     [31:0] n2100;
wire     [31:0] n2101;
wire     [31:0] n2102;
wire     [31:0] n2103;
wire     [31:0] n2104;
wire     [31:0] n2105;
wire     [31:0] n2106;
wire     [31:0] n2107;
wire     [31:0] n2108;
wire     [31:0] n2109;
wire     [31:0] n2110;
wire            n2111;
wire     [31:0] n2112;
wire     [31:0] n2113;
wire     [31:0] n2114;
wire     [31:0] n2115;
wire     [31:0] n2116;
wire     [31:0] n2117;
wire     [31:0] n2118;
wire     [31:0] n2119;
wire     [31:0] n2120;
wire     [31:0] n2121;
wire     [31:0] n2122;
wire     [31:0] n2123;
wire     [31:0] n2124;
wire     [31:0] n2125;
wire     [31:0] n2126;
wire     [31:0] n2127;
wire     [31:0] n2128;
wire     [31:0] n2129;
wire     [31:0] n2130;
wire     [31:0] n2131;
wire     [31:0] n2132;
wire     [31:0] n2133;
wire     [31:0] n2134;
wire     [31:0] n2135;
wire     [31:0] n2136;
wire     [31:0] n2137;
wire     [31:0] n2138;
wire     [31:0] n2139;
wire     [31:0] n2140;
wire     [31:0] n2141;
wire     [31:0] n2142;
wire     [31:0] n2143;
wire     [31:0] n2144;
wire     [31:0] n2145;
wire     [31:0] n2146;
wire     [31:0] n2147;
wire     [31:0] n2148;
wire     [31:0] n2149;
wire     [31:0] n2150;
wire     [31:0] n2151;
wire     [31:0] n2152;
wire     [31:0] n2153;
wire     [31:0] n2154;
wire     [31:0] n2155;
wire     [31:0] n2156;
wire     [31:0] n2157;
wire     [31:0] n2158;
wire     [31:0] n2159;
wire     [31:0] n2160;
wire     [31:0] n2161;
wire     [31:0] n2162;
wire     [31:0] n2163;
wire     [31:0] n2164;
wire     [31:0] n2165;
wire     [31:0] n2166;
wire            n2167;
wire     [31:0] n2168;
wire     [31:0] n2169;
wire     [31:0] n2170;
wire     [31:0] n2171;
wire     [31:0] n2172;
wire     [31:0] n2173;
wire     [31:0] n2174;
wire     [31:0] n2175;
wire     [31:0] n2176;
wire     [31:0] n2177;
wire     [31:0] n2178;
wire     [31:0] n2179;
wire     [31:0] n2180;
wire     [31:0] n2181;
wire     [31:0] n2182;
wire     [31:0] n2183;
wire     [31:0] n2184;
wire     [31:0] n2185;
wire     [31:0] n2186;
wire     [31:0] n2187;
wire     [31:0] n2188;
wire     [31:0] n2189;
wire     [31:0] n2190;
wire     [31:0] n2191;
wire     [31:0] n2192;
wire     [31:0] n2193;
wire     [31:0] n2194;
wire     [31:0] n2195;
wire     [31:0] n2196;
wire     [31:0] n2197;
wire     [31:0] n2198;
wire     [31:0] n2199;
wire     [31:0] n2200;
wire     [31:0] n2201;
wire     [31:0] n2202;
wire     [31:0] n2203;
wire     [31:0] n2204;
wire     [31:0] n2205;
wire     [31:0] n2206;
wire     [31:0] n2207;
wire     [31:0] n2208;
wire     [31:0] n2209;
wire     [31:0] n2210;
wire     [31:0] n2211;
wire     [31:0] n2212;
wire     [31:0] n2213;
wire     [31:0] n2214;
wire     [31:0] n2215;
wire     [31:0] n2216;
wire     [31:0] n2217;
wire     [31:0] n2218;
wire     [31:0] n2219;
wire     [31:0] n2220;
wire     [31:0] n2221;
wire     [31:0] n2222;
wire            n2223;
wire     [31:0] n2224;
wire     [31:0] n2225;
wire     [31:0] n2226;
wire     [31:0] n2227;
wire     [31:0] n2228;
wire     [31:0] n2229;
wire     [31:0] n2230;
wire     [31:0] n2231;
wire     [31:0] n2232;
wire     [31:0] n2233;
wire     [31:0] n2234;
wire     [31:0] n2235;
wire     [31:0] n2236;
wire     [31:0] n2237;
wire     [31:0] n2238;
wire     [31:0] n2239;
wire     [31:0] n2240;
wire     [31:0] n2241;
wire     [31:0] n2242;
wire     [31:0] n2243;
wire     [31:0] n2244;
wire     [31:0] n2245;
wire     [31:0] n2246;
wire     [31:0] n2247;
wire     [31:0] n2248;
wire     [31:0] n2249;
wire     [31:0] n2250;
wire     [31:0] n2251;
wire     [31:0] n2252;
wire     [31:0] n2253;
wire     [31:0] n2254;
wire     [31:0] n2255;
wire     [31:0] n2256;
wire     [31:0] n2257;
wire     [31:0] n2258;
wire     [31:0] n2259;
wire     [31:0] n2260;
wire     [31:0] n2261;
wire     [31:0] n2262;
wire     [31:0] n2263;
wire     [31:0] n2264;
wire     [31:0] n2265;
wire     [31:0] n2266;
wire     [31:0] n2267;
wire     [31:0] n2268;
wire     [31:0] n2269;
wire     [31:0] n2270;
wire     [31:0] n2271;
wire     [31:0] n2272;
wire     [31:0] n2273;
wire     [31:0] n2274;
wire     [31:0] n2275;
wire     [31:0] n2276;
wire     [31:0] n2277;
wire     [31:0] n2278;
wire            n2279;
wire     [31:0] n2280;
wire     [31:0] n2281;
wire     [31:0] n2282;
wire     [31:0] n2283;
wire     [31:0] n2284;
wire     [31:0] n2285;
wire     [31:0] n2286;
wire     [31:0] n2287;
wire     [31:0] n2288;
wire     [31:0] n2289;
wire     [31:0] n2290;
wire     [31:0] n2291;
wire     [31:0] n2292;
wire     [31:0] n2293;
wire     [31:0] n2294;
wire     [31:0] n2295;
wire     [31:0] n2296;
wire     [31:0] n2297;
wire     [31:0] n2298;
wire     [31:0] n2299;
wire     [31:0] n2300;
wire     [31:0] n2301;
wire     [31:0] n2302;
wire     [31:0] n2303;
wire     [31:0] n2304;
wire     [31:0] n2305;
wire     [31:0] n2306;
wire     [31:0] n2307;
wire     [31:0] n2308;
wire     [31:0] n2309;
wire     [31:0] n2310;
wire     [31:0] n2311;
wire     [31:0] n2312;
wire     [31:0] n2313;
wire     [31:0] n2314;
wire     [31:0] n2315;
wire     [31:0] n2316;
wire     [31:0] n2317;
wire     [31:0] n2318;
wire     [31:0] n2319;
wire     [31:0] n2320;
wire     [31:0] n2321;
wire     [31:0] n2322;
wire     [31:0] n2323;
wire     [31:0] n2324;
wire     [31:0] n2325;
wire     [31:0] n2326;
wire     [31:0] n2327;
wire     [31:0] n2328;
wire     [31:0] n2329;
wire     [31:0] n2330;
wire     [31:0] n2331;
wire     [31:0] n2332;
wire     [31:0] n2333;
wire     [31:0] n2334;
wire            n2335;
wire     [31:0] n2336;
wire     [31:0] n2337;
wire     [31:0] n2338;
wire     [31:0] n2339;
wire     [31:0] n2340;
wire     [31:0] n2341;
wire     [31:0] n2342;
wire     [31:0] n2343;
wire     [31:0] n2344;
wire     [31:0] n2345;
wire     [31:0] n2346;
wire     [31:0] n2347;
wire     [31:0] n2348;
wire     [31:0] n2349;
wire     [31:0] n2350;
wire     [31:0] n2351;
wire     [31:0] n2352;
wire     [31:0] n2353;
wire     [31:0] n2354;
wire     [31:0] n2355;
wire     [31:0] n2356;
wire     [31:0] n2357;
wire     [31:0] n2358;
wire     [31:0] n2359;
wire     [31:0] n2360;
wire     [31:0] n2361;
wire     [31:0] n2362;
wire     [31:0] n2363;
wire     [31:0] n2364;
wire     [31:0] n2365;
wire     [31:0] n2366;
wire     [31:0] n2367;
wire     [31:0] n2368;
wire     [31:0] n2369;
wire     [31:0] n2370;
wire     [31:0] n2371;
wire     [31:0] n2372;
wire     [31:0] n2373;
wire     [31:0] n2374;
wire     [31:0] n2375;
wire     [31:0] n2376;
wire     [31:0] n2377;
wire     [31:0] n2378;
wire     [31:0] n2379;
wire     [31:0] n2380;
wire     [31:0] n2381;
wire     [31:0] n2382;
wire     [31:0] n2383;
wire     [31:0] n2384;
wire     [31:0] n2385;
wire     [31:0] n2386;
wire     [31:0] n2387;
wire     [31:0] n2388;
wire     [31:0] n2389;
wire     [31:0] n2390;
wire            n2391;
wire     [31:0] n2392;
wire     [31:0] n2393;
wire     [31:0] n2394;
wire     [31:0] n2395;
wire     [31:0] n2396;
wire     [31:0] n2397;
wire     [31:0] n2398;
wire     [31:0] n2399;
wire     [31:0] n2400;
wire     [31:0] n2401;
wire     [31:0] n2402;
wire     [31:0] n2403;
wire     [31:0] n2404;
wire     [31:0] n2405;
wire     [31:0] n2406;
wire     [31:0] n2407;
wire     [31:0] n2408;
wire     [31:0] n2409;
wire     [31:0] n2410;
wire     [31:0] n2411;
wire     [31:0] n2412;
wire     [31:0] n2413;
wire     [31:0] n2414;
wire     [31:0] n2415;
wire     [31:0] n2416;
wire     [31:0] n2417;
wire     [31:0] n2418;
wire     [31:0] n2419;
wire     [31:0] n2420;
wire     [31:0] n2421;
wire     [31:0] n2422;
wire     [31:0] n2423;
wire     [31:0] n2424;
wire     [31:0] n2425;
wire     [31:0] n2426;
wire     [31:0] n2427;
wire     [31:0] n2428;
wire     [31:0] n2429;
wire     [31:0] n2430;
wire     [31:0] n2431;
wire     [31:0] n2432;
wire     [31:0] n2433;
wire     [31:0] n2434;
wire     [31:0] n2435;
wire     [31:0] n2436;
wire     [31:0] n2437;
wire     [31:0] n2438;
wire     [31:0] n2439;
wire     [31:0] n2440;
wire     [31:0] n2441;
wire     [31:0] n2442;
wire     [31:0] n2443;
wire     [31:0] n2444;
wire     [31:0] n2445;
wire     [31:0] n2446;
wire            n2447;
wire     [31:0] n2448;
wire     [31:0] n2449;
wire     [31:0] n2450;
wire     [31:0] n2451;
wire     [31:0] n2452;
wire     [31:0] n2453;
wire     [31:0] n2454;
wire     [31:0] n2455;
wire     [31:0] n2456;
wire     [31:0] n2457;
wire     [31:0] n2458;
wire     [31:0] n2459;
wire     [31:0] n2460;
wire     [31:0] n2461;
wire     [31:0] n2462;
wire     [31:0] n2463;
wire     [31:0] n2464;
wire     [31:0] n2465;
wire     [31:0] n2466;
wire     [31:0] n2467;
wire     [31:0] n2468;
wire     [31:0] n2469;
wire     [31:0] n2470;
wire     [31:0] n2471;
wire     [31:0] n2472;
wire     [31:0] n2473;
wire     [31:0] n2474;
wire     [31:0] n2475;
wire     [31:0] n2476;
wire     [31:0] n2477;
wire     [31:0] n2478;
wire     [31:0] n2479;
wire     [31:0] n2480;
wire     [31:0] n2481;
wire     [31:0] n2482;
wire     [31:0] n2483;
wire     [31:0] n2484;
wire     [31:0] n2485;
wire     [31:0] n2486;
wire     [31:0] n2487;
wire     [31:0] n2488;
wire     [31:0] n2489;
wire     [31:0] n2490;
wire     [31:0] n2491;
wire     [31:0] n2492;
wire     [31:0] n2493;
wire     [31:0] n2494;
wire     [31:0] n2495;
wire     [31:0] n2496;
wire     [31:0] n2497;
wire     [31:0] n2498;
wire     [31:0] n2499;
wire     [31:0] n2500;
wire     [31:0] n2501;
wire     [31:0] n2502;
wire            n2503;
wire     [31:0] n2504;
wire     [31:0] n2505;
wire     [31:0] n2506;
wire     [31:0] n2507;
wire     [31:0] n2508;
wire     [31:0] n2509;
wire     [31:0] n2510;
wire     [31:0] n2511;
wire     [31:0] n2512;
wire     [31:0] n2513;
wire     [31:0] n2514;
wire     [31:0] n2515;
wire     [31:0] n2516;
wire     [31:0] n2517;
wire     [31:0] n2518;
wire     [31:0] n2519;
wire     [31:0] n2520;
wire     [31:0] n2521;
wire     [31:0] n2522;
wire     [31:0] n2523;
wire     [31:0] n2524;
wire     [31:0] n2525;
wire     [31:0] n2526;
wire     [31:0] n2527;
wire     [31:0] n2528;
wire     [31:0] n2529;
wire     [31:0] n2530;
wire     [31:0] n2531;
wire     [31:0] n2532;
wire     [31:0] n2533;
wire     [31:0] n2534;
wire     [31:0] n2535;
wire     [31:0] n2536;
wire     [31:0] n2537;
wire     [31:0] n2538;
wire     [31:0] n2539;
wire     [31:0] n2540;
wire     [31:0] n2541;
wire     [31:0] n2542;
wire     [31:0] n2543;
wire     [31:0] n2544;
wire     [31:0] n2545;
wire     [31:0] n2546;
wire     [31:0] n2547;
wire     [31:0] n2548;
wire     [31:0] n2549;
wire     [31:0] n2550;
wire     [31:0] n2551;
wire     [31:0] n2552;
wire     [31:0] n2553;
wire     [31:0] n2554;
wire     [31:0] n2555;
wire     [31:0] n2556;
wire     [31:0] n2557;
wire     [31:0] n2558;
wire            n2559;
wire     [31:0] n2560;
wire     [31:0] n2561;
wire     [31:0] n2562;
wire     [31:0] n2563;
wire     [31:0] n2564;
wire     [31:0] n2565;
wire     [31:0] n2566;
wire     [31:0] n2567;
wire     [31:0] n2568;
wire     [31:0] n2569;
wire     [31:0] n2570;
wire     [31:0] n2571;
wire     [31:0] n2572;
wire     [31:0] n2573;
wire     [31:0] n2574;
wire     [31:0] n2575;
wire     [31:0] n2576;
wire     [31:0] n2577;
wire     [31:0] n2578;
wire     [31:0] n2579;
wire     [31:0] n2580;
wire     [31:0] n2581;
wire     [31:0] n2582;
wire     [31:0] n2583;
wire     [31:0] n2584;
wire     [31:0] n2585;
wire     [31:0] n2586;
wire     [31:0] n2587;
wire     [31:0] n2588;
wire     [31:0] n2589;
wire     [31:0] n2590;
wire     [31:0] n2591;
wire     [31:0] n2592;
wire     [31:0] n2593;
wire     [31:0] n2594;
wire     [31:0] n2595;
wire     [31:0] n2596;
wire     [31:0] n2597;
wire     [31:0] n2598;
wire     [31:0] n2599;
wire     [31:0] n2600;
wire     [31:0] n2601;
wire     [31:0] n2602;
wire     [31:0] n2603;
wire     [31:0] n2604;
wire     [31:0] n2605;
wire     [31:0] n2606;
wire     [31:0] n2607;
wire     [31:0] n2608;
wire     [31:0] n2609;
wire     [31:0] n2610;
wire     [31:0] n2611;
wire     [31:0] n2612;
wire     [31:0] n2613;
wire     [31:0] n2614;
wire            n2615;
wire     [31:0] n2616;
wire     [31:0] n2617;
wire     [31:0] n2618;
wire     [31:0] n2619;
wire     [31:0] n2620;
wire     [31:0] n2621;
wire     [31:0] n2622;
wire     [31:0] n2623;
wire     [31:0] n2624;
wire     [31:0] n2625;
wire     [31:0] n2626;
wire     [31:0] n2627;
wire     [31:0] n2628;
wire     [31:0] n2629;
wire     [31:0] n2630;
wire     [31:0] n2631;
wire     [31:0] n2632;
wire     [31:0] n2633;
wire     [31:0] n2634;
wire     [31:0] n2635;
wire     [31:0] n2636;
wire     [31:0] n2637;
wire     [31:0] n2638;
wire     [31:0] n2639;
wire     [31:0] n2640;
wire     [31:0] n2641;
wire     [31:0] n2642;
wire     [31:0] n2643;
wire     [31:0] n2644;
wire     [31:0] n2645;
wire     [31:0] n2646;
wire     [31:0] n2647;
wire     [31:0] n2648;
wire     [31:0] n2649;
wire     [31:0] n2650;
wire     [31:0] n2651;
wire     [31:0] n2652;
wire     [31:0] n2653;
wire     [31:0] n2654;
wire     [31:0] n2655;
wire     [31:0] n2656;
wire     [31:0] n2657;
wire     [31:0] n2658;
wire     [31:0] n2659;
wire     [31:0] n2660;
wire     [31:0] n2661;
wire     [31:0] n2662;
wire     [31:0] n2663;
wire     [31:0] n2664;
wire     [31:0] n2665;
wire     [31:0] n2666;
wire     [31:0] n2667;
wire     [31:0] n2668;
wire     [31:0] n2669;
wire     [31:0] n2670;
wire     [31:0] n2671;
wire            n2672;
wire     [31:0] n2673;
wire     [31:0] n2674;
wire     [31:0] n2675;
wire     [31:0] n2676;
wire     [31:0] n2677;
wire     [31:0] n2678;
wire     [31:0] n2679;
wire     [31:0] n2680;
wire     [31:0] n2681;
wire     [31:0] n2682;
wire     [31:0] n2683;
wire     [31:0] n2684;
wire     [31:0] n2685;
wire     [31:0] n2686;
wire     [31:0] n2687;
wire     [31:0] n2688;
wire     [31:0] n2689;
wire     [31:0] n2690;
wire     [31:0] n2691;
wire     [31:0] n2692;
wire     [31:0] n2693;
wire     [31:0] n2694;
wire     [31:0] n2695;
wire     [31:0] n2696;
wire     [31:0] n2697;
wire     [31:0] n2698;
wire     [31:0] n2699;
wire     [31:0] n2700;
wire     [31:0] n2701;
wire     [31:0] n2702;
wire     [31:0] n2703;
wire     [31:0] n2704;
wire     [31:0] n2705;
wire     [31:0] n2706;
wire     [31:0] n2707;
wire     [31:0] n2708;
wire     [31:0] n2709;
wire     [31:0] n2710;
wire     [31:0] n2711;
wire     [31:0] n2712;
wire     [31:0] n2713;
wire     [31:0] n2714;
wire     [31:0] n2715;
wire     [31:0] n2716;
wire     [31:0] n2717;
wire     [31:0] n2718;
wire     [31:0] n2719;
wire     [31:0] n2720;
wire     [31:0] n2721;
wire     [31:0] n2722;
wire     [31:0] n2723;
wire     [31:0] n2724;
wire     [31:0] n2725;
wire     [31:0] n2726;
wire     [31:0] n2727;
wire            n2728;
wire     [31:0] n2729;
wire     [31:0] n2730;
wire     [31:0] n2731;
wire     [31:0] n2732;
wire     [31:0] n2733;
wire     [31:0] n2734;
wire     [31:0] n2735;
wire     [31:0] n2736;
wire     [31:0] n2737;
wire     [31:0] n2738;
wire     [31:0] n2739;
wire     [31:0] n2740;
wire     [31:0] n2741;
wire     [31:0] n2742;
wire     [31:0] n2743;
wire     [31:0] n2744;
wire     [31:0] n2745;
wire     [31:0] n2746;
wire     [31:0] n2747;
wire     [31:0] n2748;
wire     [31:0] n2749;
wire     [31:0] n2750;
wire     [31:0] n2751;
wire     [31:0] n2752;
wire     [31:0] n2753;
wire     [31:0] n2754;
wire     [31:0] n2755;
wire     [31:0] n2756;
wire     [31:0] n2757;
wire     [31:0] n2758;
wire     [31:0] n2759;
wire     [31:0] n2760;
wire     [31:0] n2761;
wire     [31:0] n2762;
wire     [31:0] n2763;
wire     [31:0] n2764;
wire     [31:0] n2765;
wire     [31:0] n2766;
wire     [31:0] n2767;
wire     [31:0] n2768;
wire     [31:0] n2769;
wire     [31:0] n2770;
wire     [31:0] n2771;
wire     [31:0] n2772;
wire     [31:0] n2773;
wire     [31:0] n2774;
wire     [31:0] n2775;
wire     [31:0] n2776;
wire     [31:0] n2777;
wire     [31:0] n2778;
wire     [31:0] n2779;
wire     [31:0] n2780;
wire     [31:0] n2781;
wire     [31:0] n2782;
wire     [31:0] n2783;
wire            n2784;
wire     [31:0] n2785;
wire     [31:0] n2786;
wire     [31:0] n2787;
wire     [31:0] n2788;
wire     [31:0] n2789;
wire     [31:0] n2790;
wire     [31:0] n2791;
wire     [31:0] n2792;
wire     [31:0] n2793;
wire     [31:0] n2794;
wire     [31:0] n2795;
wire     [31:0] n2796;
wire     [31:0] n2797;
wire     [31:0] n2798;
wire     [31:0] n2799;
wire     [31:0] n2800;
wire     [31:0] n2801;
wire     [31:0] n2802;
wire     [31:0] n2803;
wire     [31:0] n2804;
wire     [31:0] n2805;
wire     [31:0] n2806;
wire     [31:0] n2807;
wire     [31:0] n2808;
wire     [31:0] n2809;
wire     [31:0] n2810;
wire     [31:0] n2811;
wire     [31:0] n2812;
wire     [31:0] n2813;
wire     [31:0] n2814;
wire     [31:0] n2815;
wire     [31:0] n2816;
wire     [31:0] n2817;
wire     [31:0] n2818;
wire     [31:0] n2819;
wire     [31:0] n2820;
wire     [31:0] n2821;
wire     [31:0] n2822;
wire     [31:0] n2823;
wire     [31:0] n2824;
wire     [31:0] n2825;
wire     [31:0] n2826;
wire     [31:0] n2827;
wire     [31:0] n2828;
wire     [31:0] n2829;
wire     [31:0] n2830;
wire     [31:0] n2831;
wire     [31:0] n2832;
wire     [31:0] n2833;
wire     [31:0] n2834;
wire     [31:0] n2835;
wire     [31:0] n2836;
wire     [31:0] n2837;
wire     [31:0] n2838;
wire     [31:0] n2839;
wire     [31:0] mem_addr0;
wire     [31:0] mem_data0;
wire            mem_wen0;
wire            n2840;
wire            n2841;
wire            n2842;
wire            n2843;
wire            n2844;
wire            n2845;
wire            n2846;
wire            n2847;
wire            n2848;
wire     [11:0] n2849;
wire     [31:0] n2850;
wire     [31:0] n2851;
wire     [29:0] n2852;
wire     [31:0] n2853;
wire     [31:0] n2854;
wire      [1:0] n2855;
wire     [31:0] n2856;
wire     [31:0] n2857;
wire     [31:0] n2858;
wire     [31:0] n2859;
wire     [31:0] n2860;
wire     [31:0] n2863;
wire     [31:0] n2864;
wire     [31:0] n2865;
wire            n2866;
wire     [31:0] n2867;
wire     [31:0] n2868;
wire     [31:0] n2869;
wire     [31:0] n2870;
wire     [31:0] n2871;
wire     [31:0] n2872;
wire            n2873;
wire     [31:0] n2874;
wire     [31:0] n2875;
wire     [31:0] n2876;
wire     [31:0] n2877;
wire     [31:0] n2878;
wire     [31:0] n2879;
wire clk;
wire rst;
wire step;
assign n0 =  ( Priv ) == ( 2'd1 )  ;
assign n1 = mstatus[1:1] ;
assign n2 =  ( n1 ) == ( 1'd1 )  ;
assign n3 =  ( n0 ) & ( n2 )  ;
assign n4 =  ( Priv ) < ( 2'd1 )  ;
assign n5 =  ( n3 ) | ( n4 )  ;
assign n6 =  { ( ssInt ) , ( 1'd0 ) }  ;
assign n7 =  { ( 1'd0 ) , ( n6 ) }  ;
assign n8 =  { ( msInt ) , ( n7 ) }  ;
assign n9 =  { ( 1'd0 ) , ( n8 ) }  ;
assign n10 =  { ( stInt ) , ( n9 ) }  ;
assign n11 =  { ( 1'd0 ) , ( n10 ) }  ;
assign n12 =  { ( mtInt ) , ( n11 ) }  ;
assign n13 =  { ( 1'd0 ) , ( n12 ) }  ;
assign n14 =  { ( seInt ) , ( n13 ) }  ;
assign n15 =  { ( 1'd0 ) , ( n14 ) }  ;
assign n16 =  { ( meInt ) , ( n15 ) }  ;
assign n17 =  {20'd0 , n16}  ;
assign n18 =  ( n17 ) & ( mie )  ;
assign n19 = n18[1:1] ;
assign n20 = mideleg[1:1] ;
assign n21 =  ( n19 ) & ( n20 )  ;
assign n22 =  ( n21 ) == ( 1'd1 )  ;
assign n23 =  ( n5 ) & ( n22 )  ;
assign n24 =  ( 32'd1 ) << ( 32'd1 )  ;
assign n25 =  ( Priv ) == ( 2'd3 )  ;
assign n26 = mstatus[3:3] ;
assign n27 =  ( n26 ) == ( 1'd1 )  ;
assign n28 =  ( n25 ) & ( n27 )  ;
assign n29 =  ( Priv ) < ( 2'd3 )  ;
assign n30 =  ( n28 ) | ( n29 )  ;
assign n31 = ~ ( n20 ) ;
assign n32 =  ( n19 ) & ( n31 )  ;
assign n33 =  ( n32 ) == ( 1'd1 )  ;
assign n34 =  ( n30 ) & ( n33 )  ;
assign n35 = n18[3:3] ;
assign n36 = mideleg[3:3] ;
assign n37 = ~ ( n36 ) ;
assign n38 =  ( n35 ) & ( n37 )  ;
assign n39 =  ( n38 ) == ( 1'd1 )  ;
assign n40 =  ( n30 ) & ( n39 )  ;
assign n41 =  ( 32'd1 ) << ( 32'd3 )  ;
assign n42 = n18[5:5] ;
assign n43 = mideleg[5:5] ;
assign n44 =  ( n42 ) & ( n43 )  ;
assign n45 =  ( n44 ) == ( 1'd1 )  ;
assign n46 =  ( n5 ) & ( n45 )  ;
assign n47 =  ( 32'd1 ) << ( 32'd5 )  ;
assign n48 = ~ ( n43 ) ;
assign n49 =  ( n42 ) & ( n48 )  ;
assign n50 =  ( n49 ) == ( 1'd1 )  ;
assign n51 =  ( n30 ) & ( n50 )  ;
assign n52 = n18[7:7] ;
assign n53 = mideleg[7:7] ;
assign n54 = ~ ( n53 ) ;
assign n55 =  ( n52 ) & ( n54 )  ;
assign n56 =  ( n55 ) == ( 1'd1 )  ;
assign n57 =  ( n30 ) & ( n56 )  ;
assign n58 =  ( 32'd1 ) << ( 32'd7 )  ;
assign n59 = n18[9:9] ;
assign n60 = mideleg[9:9] ;
assign n61 =  ( n59 ) & ( n60 )  ;
assign n62 =  ( n61 ) == ( 1'd1 )  ;
assign n63 =  ( n5 ) & ( n62 )  ;
assign n64 =  ( 32'd1 ) << ( 32'd9 )  ;
assign n65 = ~ ( n60 ) ;
assign n66 =  ( n59 ) & ( n65 )  ;
assign n67 =  ( n66 ) == ( 1'd1 )  ;
assign n68 =  ( n30 ) & ( n67 )  ;
assign n69 = n18[11:11] ;
assign n70 = mideleg[11:11] ;
assign n71 = ~ ( n70 ) ;
assign n72 =  ( n69 ) & ( n71 )  ;
assign n73 =  ( n72 ) == ( 1'd1 )  ;
assign n74 =  ( n30 ) & ( n73 )  ;
assign n75 =  ( 32'd1 ) << ( 32'd11 )  ;
assign n76 =  ( n74 ) ? ( n75 ) : ( 32'd0 ) ;
assign n77 =  ( n68 ) ? ( n64 ) : ( n76 ) ;
assign n78 =  ( n63 ) ? ( n64 ) : ( n77 ) ;
assign n79 =  ( n57 ) ? ( n58 ) : ( n78 ) ;
assign n80 =  ( n51 ) ? ( n47 ) : ( n79 ) ;
assign n81 =  ( n46 ) ? ( n47 ) : ( n80 ) ;
assign n82 =  ( n40 ) ? ( n41 ) : ( n81 ) ;
assign n83 =  ( n34 ) ? ( n24 ) : ( n82 ) ;
assign n84__int_trap_select =  ( n23 ) ? ( n24 ) : ( n83 ) ;
assign n85 = n84__int_trap_select[1:1] ;
assign n86 =  ( n85 ) & ( n20 )  ;
assign n87 = n84__int_trap_select[5:5] ;
assign n88 =  ( n87 ) & ( n43 )  ;
assign n89 =  ( n86 ) | ( n88 )  ;
assign n90 = n84__int_trap_select[9:9] ;
assign n91 =  ( n90 ) & ( n60 )  ;
assign n92 =  ( n89 ) | ( n91 )  ;
assign n93 =  ( n92 ) == ( 1'd1 )  ;
assign n94 = n84__int_trap_select[3:3] ;
assign n95 = n84__int_trap_select[7:7] ;
assign n96 =  ( n94 ) | ( n95 )  ;
assign n97 = n84__int_trap_select[11:11] ;
assign n98 =  ( n96 ) | ( n97 )  ;
assign n99 =  ( n85 ) & ( n31 )  ;
assign n100 =  ( n87 ) & ( n48 )  ;
assign n101 =  ( n99 ) | ( n100 )  ;
assign n102 =  ( n90 ) & ( n65 )  ;
assign n103 =  ( n101 ) | ( n102 )  ;
assign n104 =  ( n98 ) | ( n103 )  ;
assign n105 =  ( n104 ) == ( 1'd1 )  ;
assign n106__take_int_sig =  ( n93 ) | ( n105 )  ;
assign n107 = pc[1:0] ;
assign n108 =  ( n107 ) != ( 2'd0 )  ;
assign n109 = pc[31:2] ;
assign n110 =  {2'd0 , n109}  ;
assign mem_addr_n111 = n110 ;
assign n113 = mem_data_n112 ;
assign n114 =  ( n113 ) == ( 32'd270532723 )  ;
assign n115 =  ( n113 ) == ( 32'd807403635 )  ;
assign n116 =  ( n114 ) | ( n115 )  ;
assign n117 = mepc[1:0] ;
assign n118 =  ( n117 ) != ( 2'd0 )  ;
assign n119 =  ( n115 ) & ( n118 )  ;
assign n120 = sepc[1:0] ;
assign n121 =  ( n120 ) != ( 2'd0 )  ;
assign n122 =  ( n114 ) & ( n121 )  ;
assign n123 =  ( n119 ) | ( n122 )  ;
assign n124 =  ( n116 ) & ( n123 )  ;
assign n125 =  ( n108 ) | ( n124 )  ;
assign n126 =  ( 32'd57347 ) & ( n113 )  ;
assign n127 =  ( 32'd57346 ) == ( n126 )  ;
assign n128 =  ( 32'd49154 ) == ( n126 )  ;
assign n129 =  ( 32'd40962 ) == ( n126 )  ;
assign n130 =  ( 32'd61443 ) & ( n113 )  ;
assign n131 =  ( 32'd36866 ) == ( n130 )  ;
assign n132 =  ( 32'd32770 ) == ( n130 )  ;
assign n133 =  ( 32'd24578 ) == ( n126 )  ;
assign n134 =  ( 32'd16386 ) == ( n126 )  ;
assign n135 =  ( 32'd8194 ) == ( n126 )  ;
assign n136 =  ( 32'd2 ) == ( n126 )  ;
assign n137 =  ( 32'd57345 ) == ( n126 )  ;
assign n138 =  ( 32'd49153 ) == ( n126 )  ;
assign n139 =  ( 32'd40961 ) == ( n126 )  ;
assign n140 =  ( 32'd64611 ) & ( n113 )  ;
assign n141 =  ( 32'd39969 ) == ( n140 )  ;
assign n142 =  ( 32'd39937 ) == ( n140 )  ;
assign n143 =  ( 32'd35937 ) == ( n140 )  ;
assign n144 =  ( 32'd35905 ) == ( n140 )  ;
assign n145 =  ( 32'd35873 ) == ( n140 )  ;
assign n146 =  ( 32'd35841 ) == ( n140 )  ;
assign n147 =  ( 32'd60419 ) & ( n113 )  ;
assign n148 =  ( 32'd34817 ) == ( n147 )  ;
assign n149 =  ( 32'd33793 ) == ( n147 )  ;
assign n150 =  ( 32'd32769 ) == ( n147 )  ;
assign n151 =  ( 32'd24577 ) == ( n126 )  ;
assign n152 =  ( 32'd16385 ) == ( n126 )  ;
assign n153 =  ( 32'd8193 ) == ( n126 )  ;
assign n154 =  ( 32'd1 ) == ( n126 )  ;
assign n155 =  ( 32'd57344 ) == ( n126 )  ;
assign n156 =  ( 32'd49152 ) == ( n126 )  ;
assign n157 =  ( 32'd40960 ) == ( n126 )  ;
assign n158 =  ( 32'd24576 ) == ( n126 )  ;
assign n159 =  ( 32'd16384 ) == ( n126 )  ;
assign n160 =  ( 32'd8192 ) == ( n126 )  ;
assign n161 =  ( 32'd0 ) == ( n126 )  ;
assign n162 =  ( 32'd65535 ) & ( n113 )  ;
assign n163 =  ( 32'd36866 ) == ( n162 )  ;
assign n164 =  ( 32'd61567 ) & ( n113 )  ;
assign n165 =  ( 32'd36866 ) == ( n164 )  ;
assign n166 =  ( 32'd32770 ) == ( n164 )  ;
assign n167 =  ( 32'd61315 ) & ( n113 )  ;
assign n168 =  ( 32'd24833 ) == ( n167 )  ;
assign n169 =  ( 32'd1 ) == ( n162 )  ;
assign n170 =  ( 32'd100663423 ) & ( n113 )  ;
assign n171 =  ( 32'd33554511 ) == ( n170 )  ;
assign n172 =  ( 32'd33554507 ) == ( n170 )  ;
assign n173 =  ( 32'd33554503 ) == ( n170 )  ;
assign n174 =  ( 32'd33554499 ) == ( n170 )  ;
assign n175 =  ( 32'd79 ) == ( n170 )  ;
assign n176 =  ( 32'd75 ) == ( n170 )  ;
assign n177 =  ( 32'd71 ) == ( n170 )  ;
assign n178 =  ( 32'd67 ) == ( n170 )  ;
assign n179 =  ( 32'd28799 ) & ( n113 )  ;
assign n180 =  ( 32'd12327 ) == ( n179 )  ;
assign n181 =  ( 32'd8231 ) == ( n179 )  ;
assign n182 =  ( 32'd12295 ) == ( n179 )  ;
assign n183 =  ( 32'd8199 ) == ( n179 )  ;
assign n184 =  ( 32'd4293947519 ) & ( n113 )  ;
assign n185 =  ( 32'd4060086355 ) == ( n184 )  ;
assign n186 =  ( 32'd4293918847 ) & ( n113 )  ;
assign n187 =  ( 32'd3526361171 ) == ( n186 )  ;
assign n188 =  ( 32'd3525312595 ) == ( n186 )  ;
assign n189 =  ( 32'd3524264019 ) == ( n186 )  ;
assign n190 =  ( 32'd3523215443 ) == ( n186 )  ;
assign n191 =  ( 32'd4026531923 ) == ( n184 )  ;
assign n192 =  ( 32'd3492806739 ) == ( n186 )  ;
assign n193 =  ( 32'd3491758163 ) == ( n186 )  ;
assign n194 =  ( 32'd3490709587 ) == ( n186 )  ;
assign n195 =  ( 32'd3489661011 ) == ( n186 )  ;
assign n196 =  ( 32'd3791654995 ) == ( n184 )  ;
assign n197 =  ( 32'd3791650899 ) == ( n184 )  ;
assign n198 =  ( 32'd3257925715 ) == ( n186 )  ;
assign n199 =  ( 32'd3256877139 ) == ( n186 )  ;
assign n200 =  ( 32'd3255828563 ) == ( n186 )  ;
assign n201 =  ( 32'd3254779987 ) == ( n186 )  ;
assign n202 =  ( 32'd3758100563 ) == ( n184 )  ;
assign n203 =  ( 32'd3758096467 ) == ( n184 )  ;
assign n204 =  ( 32'd3224371283 ) == ( n186 )  ;
assign n205 =  ( 32'd3223322707 ) == ( n186 )  ;
assign n206 =  ( 32'd3222274131 ) == ( n186 )  ;
assign n207 =  ( 32'd3221225555 ) == ( n186 )  ;
assign n208 =  ( 32'd4261441663 ) & ( n113 )  ;
assign n209 =  ( 32'd2717917267 ) == ( n208 )  ;
assign n210 =  ( 32'd2717913171 ) == ( n208 )  ;
assign n211 =  ( 32'd2717909075 ) == ( n208 )  ;
assign n212 =  ( 32'd2684362835 ) == ( n208 )  ;
assign n213 =  ( 32'd2684358739 ) == ( n208 )  ;
assign n214 =  ( 32'd2684354643 ) == ( n208 )  ;
assign n215 =  ( 32'd1509949523 ) == ( n186 )  ;
assign n216 =  ( 32'd1107296339 ) == ( n186 )  ;
assign n217 =  ( 32'd1074790483 ) == ( n186 )  ;
assign n218 =  ( 32'd704647251 ) == ( n208 )  ;
assign n219 =  ( 32'd704643155 ) == ( n208 )  ;
assign n220 =  ( 32'd570433619 ) == ( n208 )  ;
assign n221 =  ( 32'd570429523 ) == ( n208 )  ;
assign n222 =  ( 32'd570425427 ) == ( n208 )  ;
assign n223 =  ( 32'd4261412991 ) & ( n113 )  ;
assign n224 =  ( 32'd436207699 ) == ( n223 )  ;
assign n225 =  ( 32'd301989971 ) == ( n223 )  ;
assign n226 =  ( 32'd167772243 ) == ( n223 )  ;
assign n227 =  ( 32'd33554515 ) == ( n223 )  ;
assign n228 =  ( 32'd1476395091 ) == ( n186 )  ;
assign n229 =  ( 32'd671092819 ) == ( n208 )  ;
assign n230 =  ( 32'd671088723 ) == ( n208 )  ;
assign n231 =  ( 32'd536879187 ) == ( n208 )  ;
assign n232 =  ( 32'd536875091 ) == ( n208 )  ;
assign n233 =  ( 32'd536870995 ) == ( n208 )  ;
assign n234 =  ( 32'd402653267 ) == ( n223 )  ;
assign n235 =  ( 32'd268435539 ) == ( n223 )  ;
assign n236 =  ( 32'd134217811 ) == ( n223 )  ;
assign n237 =  ( 32'd83 ) == ( n223 )  ;
assign n238 =  ( 32'd28787 ) == ( n179 )  ;
assign n239 =  ( 32'd24691 ) == ( n179 )  ;
assign n240 =  ( 32'd20595 ) == ( n179 )  ;
assign n241 =  ( 32'd12403 ) == ( n179 )  ;
assign n242 =  ( 32'd8307 ) == ( n179 )  ;
assign n243 =  ( 32'd4211 ) == ( n179 )  ;
assign n244 =  ( 32'd4294967295 ) & ( n113 )  ;
assign n245 =  ( 32'd273678451 ) == ( n244 )  ;
assign n246 =  ( 32'd4293951487 ) & ( n113 )  ;
assign n247 =  ( 32'd272629875 ) == ( n246 )  ;
assign n248 =  ( 32'd2065694835 ) == ( n244 )  ;
assign n249 =  ( 32'd807403635 ) == ( n244 )  ;
assign n250 =  ( 32'd538968179 ) == ( n244 )  ;
assign n251 =  ( 32'd270532723 ) == ( n244 )  ;
assign n252 =  ( 32'd2097267 ) == ( n244 )  ;
assign n253 =  ( 32'd1048691 ) == ( n244 )  ;
assign n254 =  ( 32'd115 ) == ( n244 )  ;
assign n255 =  ( 32'd4160778367 ) & ( n113 )  ;
assign n256 =  ( 32'd402665519 ) == ( n255 )  ;
assign n257 =  ( 32'd4193284223 ) & ( n113 )  ;
assign n258 =  ( 32'd268447791 ) == ( n257 )  ;
assign n259 =  ( 32'd134230063 ) == ( n255 )  ;
assign n260 =  ( 32'd3758108719 ) == ( n255 )  ;
assign n261 =  ( 32'd3221237807 ) == ( n255 )  ;
assign n262 =  ( 32'd2684366895 ) == ( n255 )  ;
assign n263 =  ( 32'd2147495983 ) == ( n255 )  ;
assign n264 =  ( 32'd1610625071 ) == ( n255 )  ;
assign n265 =  ( 32'd1073754159 ) == ( n255 )  ;
assign n266 =  ( 32'd536883247 ) == ( n255 )  ;
assign n267 =  ( 32'd12335 ) == ( n255 )  ;
assign n268 =  ( 32'd402661423 ) == ( n255 )  ;
assign n269 =  ( 32'd268443695 ) == ( n257 )  ;
assign n270 =  ( 32'd134225967 ) == ( n255 )  ;
assign n271 =  ( 32'd3758104623 ) == ( n255 )  ;
assign n272 =  ( 32'd3221233711 ) == ( n255 )  ;
assign n273 =  ( 32'd2684362799 ) == ( n255 )  ;
assign n274 =  ( 32'd2147491887 ) == ( n255 )  ;
assign n275 =  ( 32'd1610620975 ) == ( n255 )  ;
assign n276 =  ( 32'd1073750063 ) == ( n255 )  ;
assign n277 =  ( 32'd536879151 ) == ( n255 )  ;
assign n278 =  ( 32'd8239 ) == ( n255 )  ;
assign n279 =  ( 32'd33583163 ) == ( n208 )  ;
assign n280 =  ( 32'd33579067 ) == ( n208 )  ;
assign n281 =  ( 32'd33574971 ) == ( n208 )  ;
assign n282 =  ( 32'd33570875 ) == ( n208 )  ;
assign n283 =  ( 32'd33554491 ) == ( n208 )  ;
assign n284 =  ( 32'd33583155 ) == ( n208 )  ;
assign n285 =  ( 32'd33579059 ) == ( n208 )  ;
assign n286 =  ( 32'd33574963 ) == ( n208 )  ;
assign n287 =  ( 32'd33570867 ) == ( n208 )  ;
assign n288 =  ( 32'd33566771 ) == ( n208 )  ;
assign n289 =  ( 32'd33562675 ) == ( n208 )  ;
assign n290 =  ( 32'd33558579 ) == ( n208 )  ;
assign n291 =  ( 32'd33554483 ) == ( n208 )  ;
assign n292 =  ( 32'd4111 ) == ( n179 )  ;
assign n293 =  ( 32'd15 ) == ( n179 )  ;
assign n294 =  ( 32'd12323 ) == ( n179 )  ;
assign n295 =  ( 32'd8227 ) == ( n179 )  ;
assign n296 =  ( 32'd4131 ) == ( n179 )  ;
assign n297 =  ( 32'd35 ) == ( n179 )  ;
assign n298 =  ( 32'd24579 ) == ( n179 )  ;
assign n299 =  ( 32'd20483 ) == ( n179 )  ;
assign n300 =  ( 32'd16387 ) == ( n179 )  ;
assign n301 =  ( 32'd12291 ) == ( n179 )  ;
assign n302 =  ( 32'd8195 ) == ( n179 )  ;
assign n303 =  ( 32'd4099 ) == ( n179 )  ;
assign n304 =  ( 32'd3 ) == ( n179 )  ;
assign n305 =  ( 32'd1073762363 ) == ( n208 )  ;
assign n306 =  ( 32'd20539 ) == ( n208 )  ;
assign n307 =  ( 32'd4155 ) == ( n208 )  ;
assign n308 =  ( 32'd1073741883 ) == ( n208 )  ;
assign n309 =  ( 32'd59 ) == ( n208 )  ;
assign n310 =  ( 32'd1073762331 ) == ( n208 )  ;
assign n311 =  ( 32'd20507 ) == ( n208 )  ;
assign n312 =  ( 32'd4123 ) == ( n208 )  ;
assign n313 =  ( 32'd27 ) == ( n179 )  ;
assign n314 =  ( 32'd28723 ) == ( n208 )  ;
assign n315 =  ( 32'd24627 ) == ( n208 )  ;
assign n316 =  ( 32'd1073762355 ) == ( n208 )  ;
assign n317 =  ( 32'd20531 ) == ( n208 )  ;
assign n318 =  ( 32'd16435 ) == ( n208 )  ;
assign n319 =  ( 32'd12339 ) == ( n208 )  ;
assign n320 =  ( 32'd8243 ) == ( n208 )  ;
assign n321 =  ( 32'd4147 ) == ( n208 )  ;
assign n322 =  ( 32'd1073741875 ) == ( n208 )  ;
assign n323 =  ( 32'd51 ) == ( n208 )  ;
assign n324 =  ( 32'd28691 ) == ( n179 )  ;
assign n325 =  ( 32'd24595 ) == ( n179 )  ;
assign n326 =  ( 32'd4227887231 ) & ( n113 )  ;
assign n327 =  ( 32'd1073762323 ) == ( n326 )  ;
assign n328 =  ( 32'd20499 ) == ( n326 )  ;
assign n329 =  ( 32'd16403 ) == ( n179 )  ;
assign n330 =  ( 32'd12307 ) == ( n179 )  ;
assign n331 =  ( 32'd8211 ) == ( n179 )  ;
assign n332 =  ( 32'd4115 ) == ( n326 )  ;
assign n333 =  ( 32'd19 ) == ( n179 )  ;
assign n334 =  ( 32'd127 ) & ( n113 )  ;
assign n335 =  ( 32'd23 ) == ( n334 )  ;
assign n336 =  ( 32'd55 ) == ( n334 )  ;
assign n337 =  ( 32'd111 ) == ( n334 )  ;
assign n338 =  ( 32'd103 ) == ( n179 )  ;
assign n339 =  ( 32'd28771 ) == ( n179 )  ;
assign n340 =  ( 32'd24675 ) == ( n179 )  ;
assign n341 =  ( 32'd20579 ) == ( n179 )  ;
assign n342 =  ( 32'd16483 ) == ( n179 )  ;
assign n343 =  ( 32'd4195 ) == ( n179 )  ;
assign n344 =  ( 32'd99 ) == ( n179 )  ;
assign n345 =  ( n344 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n346 =  ( n343 ) ? ( 1'd0 ) : ( n345 ) ;
assign n347 =  ( n342 ) ? ( 1'd0 ) : ( n346 ) ;
assign n348 =  ( n341 ) ? ( 1'd0 ) : ( n347 ) ;
assign n349 =  ( n340 ) ? ( 1'd0 ) : ( n348 ) ;
assign n350 =  ( n339 ) ? ( 1'd0 ) : ( n349 ) ;
assign n351 =  ( n338 ) ? ( 1'd0 ) : ( n350 ) ;
assign n352 =  ( n337 ) ? ( 1'd0 ) : ( n351 ) ;
assign n353 =  ( n336 ) ? ( 1'd0 ) : ( n352 ) ;
assign n354 =  ( n335 ) ? ( 1'd0 ) : ( n353 ) ;
assign n355 =  ( n333 ) ? ( 1'd0 ) : ( n354 ) ;
assign n356 =  ( n332 ) ? ( 1'd0 ) : ( n355 ) ;
assign n357 =  ( n331 ) ? ( 1'd0 ) : ( n356 ) ;
assign n358 =  ( n330 ) ? ( 1'd0 ) : ( n357 ) ;
assign n359 =  ( n329 ) ? ( 1'd0 ) : ( n358 ) ;
assign n360 =  ( n328 ) ? ( 1'd0 ) : ( n359 ) ;
assign n361 =  ( n327 ) ? ( 1'd0 ) : ( n360 ) ;
assign n362 =  ( n325 ) ? ( 1'd0 ) : ( n361 ) ;
assign n363 =  ( n324 ) ? ( 1'd0 ) : ( n362 ) ;
assign n364 =  ( n323 ) ? ( 1'd0 ) : ( n363 ) ;
assign n365 =  ( n322 ) ? ( 1'd0 ) : ( n364 ) ;
assign n366 =  ( n321 ) ? ( 1'd0 ) : ( n365 ) ;
assign n367 =  ( n320 ) ? ( 1'd0 ) : ( n366 ) ;
assign n368 =  ( n319 ) ? ( 1'd0 ) : ( n367 ) ;
assign n369 =  ( n318 ) ? ( 1'd0 ) : ( n368 ) ;
assign n370 =  ( n317 ) ? ( 1'd0 ) : ( n369 ) ;
assign n371 =  ( n316 ) ? ( 1'd0 ) : ( n370 ) ;
assign n372 =  ( n315 ) ? ( 1'd0 ) : ( n371 ) ;
assign n373 =  ( n314 ) ? ( 1'd0 ) : ( n372 ) ;
assign n374 =  ( n313 ) ? ( 1'd0 ) : ( n373 ) ;
assign n375 =  ( n312 ) ? ( 1'd0 ) : ( n374 ) ;
assign n376 =  ( n311 ) ? ( 1'd0 ) : ( n375 ) ;
assign n377 =  ( n310 ) ? ( 1'd0 ) : ( n376 ) ;
assign n378 =  ( n309 ) ? ( 1'd0 ) : ( n377 ) ;
assign n379 =  ( n308 ) ? ( 1'd0 ) : ( n378 ) ;
assign n380 =  ( n307 ) ? ( 1'd0 ) : ( n379 ) ;
assign n381 =  ( n306 ) ? ( 1'd0 ) : ( n380 ) ;
assign n382 =  ( n305 ) ? ( 1'd0 ) : ( n381 ) ;
assign n383 =  ( n304 ) ? ( 1'd0 ) : ( n382 ) ;
assign n384 =  ( n303 ) ? ( 1'd0 ) : ( n383 ) ;
assign n385 =  ( n302 ) ? ( 1'd0 ) : ( n384 ) ;
assign n386 =  ( n301 ) ? ( 1'd0 ) : ( n385 ) ;
assign n387 =  ( n300 ) ? ( 1'd0 ) : ( n386 ) ;
assign n388 =  ( n299 ) ? ( 1'd0 ) : ( n387 ) ;
assign n389 =  ( n298 ) ? ( 1'd0 ) : ( n388 ) ;
assign n390 =  ( n297 ) ? ( 1'd0 ) : ( n389 ) ;
assign n391 =  ( n296 ) ? ( 1'd0 ) : ( n390 ) ;
assign n392 =  ( n295 ) ? ( 1'd0 ) : ( n391 ) ;
assign n393 =  ( n294 ) ? ( 1'd0 ) : ( n392 ) ;
assign n394 =  ( n293 ) ? ( 1'd0 ) : ( n393 ) ;
assign n395 =  ( n292 ) ? ( 1'd0 ) : ( n394 ) ;
assign n396 =  ( n291 ) ? ( 1'd0 ) : ( n395 ) ;
assign n397 =  ( n290 ) ? ( 1'd0 ) : ( n396 ) ;
assign n398 =  ( n289 ) ? ( 1'd0 ) : ( n397 ) ;
assign n399 =  ( n288 ) ? ( 1'd0 ) : ( n398 ) ;
assign n400 =  ( n287 ) ? ( 1'd0 ) : ( n399 ) ;
assign n401 =  ( n286 ) ? ( 1'd0 ) : ( n400 ) ;
assign n402 =  ( n285 ) ? ( 1'd0 ) : ( n401 ) ;
assign n403 =  ( n284 ) ? ( 1'd0 ) : ( n402 ) ;
assign n404 =  ( n283 ) ? ( 1'd0 ) : ( n403 ) ;
assign n405 =  ( n282 ) ? ( 1'd0 ) : ( n404 ) ;
assign n406 =  ( n281 ) ? ( 1'd0 ) : ( n405 ) ;
assign n407 =  ( n280 ) ? ( 1'd0 ) : ( n406 ) ;
assign n408 =  ( n279 ) ? ( 1'd0 ) : ( n407 ) ;
assign n409 =  ( n278 ) ? ( 1'd0 ) : ( n408 ) ;
assign n410 =  ( n277 ) ? ( 1'd0 ) : ( n409 ) ;
assign n411 =  ( n276 ) ? ( 1'd0 ) : ( n410 ) ;
assign n412 =  ( n275 ) ? ( 1'd0 ) : ( n411 ) ;
assign n413 =  ( n274 ) ? ( 1'd0 ) : ( n412 ) ;
assign n414 =  ( n273 ) ? ( 1'd0 ) : ( n413 ) ;
assign n415 =  ( n272 ) ? ( 1'd0 ) : ( n414 ) ;
assign n416 =  ( n271 ) ? ( 1'd0 ) : ( n415 ) ;
assign n417 =  ( n270 ) ? ( 1'd0 ) : ( n416 ) ;
assign n418 =  ( n269 ) ? ( 1'd0 ) : ( n417 ) ;
assign n419 =  ( n268 ) ? ( 1'd0 ) : ( n418 ) ;
assign n420 =  ( n267 ) ? ( 1'd0 ) : ( n419 ) ;
assign n421 =  ( n266 ) ? ( 1'd0 ) : ( n420 ) ;
assign n422 =  ( n265 ) ? ( 1'd0 ) : ( n421 ) ;
assign n423 =  ( n264 ) ? ( 1'd0 ) : ( n422 ) ;
assign n424 =  ( n263 ) ? ( 1'd0 ) : ( n423 ) ;
assign n425 =  ( n262 ) ? ( 1'd0 ) : ( n424 ) ;
assign n426 =  ( n261 ) ? ( 1'd0 ) : ( n425 ) ;
assign n427 =  ( n260 ) ? ( 1'd0 ) : ( n426 ) ;
assign n428 =  ( n259 ) ? ( 1'd0 ) : ( n427 ) ;
assign n429 =  ( n258 ) ? ( 1'd0 ) : ( n428 ) ;
assign n430 =  ( n256 ) ? ( 1'd0 ) : ( n429 ) ;
assign n431 =  ( n254 ) ? ( 1'd0 ) : ( n430 ) ;
assign n432 =  ( n253 ) ? ( 1'd0 ) : ( n431 ) ;
assign n433 =  ( n252 ) ? ( 1'd0 ) : ( n432 ) ;
assign n434 =  ( n251 ) ? ( 1'd0 ) : ( n433 ) ;
assign n435 =  ( n250 ) ? ( 1'd0 ) : ( n434 ) ;
assign n436 =  ( n249 ) ? ( 1'd0 ) : ( n435 ) ;
assign n437 =  ( n248 ) ? ( 1'd0 ) : ( n436 ) ;
assign n438 =  ( n247 ) ? ( 1'd0 ) : ( n437 ) ;
assign n439 =  ( n245 ) ? ( 1'd0 ) : ( n438 ) ;
assign n440 =  ( n243 ) ? ( 1'd0 ) : ( n439 ) ;
assign n441 =  ( n242 ) ? ( 1'd0 ) : ( n440 ) ;
assign n442 =  ( n241 ) ? ( 1'd0 ) : ( n441 ) ;
assign n443 =  ( n240 ) ? ( 1'd0 ) : ( n442 ) ;
assign n444 =  ( n239 ) ? ( 1'd0 ) : ( n443 ) ;
assign n445 =  ( n238 ) ? ( 1'd0 ) : ( n444 ) ;
assign n446 =  ( n237 ) ? ( 1'd0 ) : ( n445 ) ;
assign n447 =  ( n236 ) ? ( 1'd0 ) : ( n446 ) ;
assign n448 =  ( n235 ) ? ( 1'd0 ) : ( n447 ) ;
assign n449 =  ( n234 ) ? ( 1'd0 ) : ( n448 ) ;
assign n450 =  ( n233 ) ? ( 1'd0 ) : ( n449 ) ;
assign n451 =  ( n232 ) ? ( 1'd0 ) : ( n450 ) ;
assign n452 =  ( n231 ) ? ( 1'd0 ) : ( n451 ) ;
assign n453 =  ( n230 ) ? ( 1'd0 ) : ( n452 ) ;
assign n454 =  ( n229 ) ? ( 1'd0 ) : ( n453 ) ;
assign n455 =  ( n228 ) ? ( 1'd0 ) : ( n454 ) ;
assign n456 =  ( n227 ) ? ( 1'd0 ) : ( n455 ) ;
assign n457 =  ( n226 ) ? ( 1'd0 ) : ( n456 ) ;
assign n458 =  ( n225 ) ? ( 1'd0 ) : ( n457 ) ;
assign n459 =  ( n224 ) ? ( 1'd0 ) : ( n458 ) ;
assign n460 =  ( n222 ) ? ( 1'd0 ) : ( n459 ) ;
assign n461 =  ( n221 ) ? ( 1'd0 ) : ( n460 ) ;
assign n462 =  ( n220 ) ? ( 1'd0 ) : ( n461 ) ;
assign n463 =  ( n219 ) ? ( 1'd0 ) : ( n462 ) ;
assign n464 =  ( n218 ) ? ( 1'd0 ) : ( n463 ) ;
assign n465 =  ( n217 ) ? ( 1'd0 ) : ( n464 ) ;
assign n466 =  ( n216 ) ? ( 1'd0 ) : ( n465 ) ;
assign n467 =  ( n215 ) ? ( 1'd0 ) : ( n466 ) ;
assign n468 =  ( n214 ) ? ( 1'd0 ) : ( n467 ) ;
assign n469 =  ( n213 ) ? ( 1'd0 ) : ( n468 ) ;
assign n470 =  ( n212 ) ? ( 1'd0 ) : ( n469 ) ;
assign n471 =  ( n211 ) ? ( 1'd0 ) : ( n470 ) ;
assign n472 =  ( n210 ) ? ( 1'd0 ) : ( n471 ) ;
assign n473 =  ( n209 ) ? ( 1'd0 ) : ( n472 ) ;
assign n474 =  ( n207 ) ? ( 1'd0 ) : ( n473 ) ;
assign n475 =  ( n206 ) ? ( 1'd0 ) : ( n474 ) ;
assign n476 =  ( n205 ) ? ( 1'd0 ) : ( n475 ) ;
assign n477 =  ( n204 ) ? ( 1'd0 ) : ( n476 ) ;
assign n478 =  ( n203 ) ? ( 1'd0 ) : ( n477 ) ;
assign n479 =  ( n202 ) ? ( 1'd0 ) : ( n478 ) ;
assign n480 =  ( n201 ) ? ( 1'd0 ) : ( n479 ) ;
assign n481 =  ( n200 ) ? ( 1'd0 ) : ( n480 ) ;
assign n482 =  ( n199 ) ? ( 1'd0 ) : ( n481 ) ;
assign n483 =  ( n198 ) ? ( 1'd0 ) : ( n482 ) ;
assign n484 =  ( n197 ) ? ( 1'd0 ) : ( n483 ) ;
assign n485 =  ( n196 ) ? ( 1'd0 ) : ( n484 ) ;
assign n486 =  ( n195 ) ? ( 1'd0 ) : ( n485 ) ;
assign n487 =  ( n194 ) ? ( 1'd0 ) : ( n486 ) ;
assign n488 =  ( n193 ) ? ( 1'd0 ) : ( n487 ) ;
assign n489 =  ( n192 ) ? ( 1'd0 ) : ( n488 ) ;
assign n490 =  ( n191 ) ? ( 1'd0 ) : ( n489 ) ;
assign n491 =  ( n190 ) ? ( 1'd0 ) : ( n490 ) ;
assign n492 =  ( n189 ) ? ( 1'd0 ) : ( n491 ) ;
assign n493 =  ( n188 ) ? ( 1'd0 ) : ( n492 ) ;
assign n494 =  ( n187 ) ? ( 1'd0 ) : ( n493 ) ;
assign n495 =  ( n185 ) ? ( 1'd0 ) : ( n494 ) ;
assign n496 =  ( n183 ) ? ( 1'd0 ) : ( n495 ) ;
assign n497 =  ( n182 ) ? ( 1'd0 ) : ( n496 ) ;
assign n498 =  ( n181 ) ? ( 1'd0 ) : ( n497 ) ;
assign n499 =  ( n180 ) ? ( 1'd0 ) : ( n498 ) ;
assign n500 =  ( n178 ) ? ( 1'd0 ) : ( n499 ) ;
assign n501 =  ( n177 ) ? ( 1'd0 ) : ( n500 ) ;
assign n502 =  ( n176 ) ? ( 1'd0 ) : ( n501 ) ;
assign n503 =  ( n175 ) ? ( 1'd0 ) : ( n502 ) ;
assign n504 =  ( n174 ) ? ( 1'd0 ) : ( n503 ) ;
assign n505 =  ( n173 ) ? ( 1'd0 ) : ( n504 ) ;
assign n506 =  ( n172 ) ? ( 1'd0 ) : ( n505 ) ;
assign n507 =  ( n171 ) ? ( 1'd0 ) : ( n506 ) ;
assign n508 =  ( n169 ) ? ( 1'd0 ) : ( n507 ) ;
assign n509 =  ( n168 ) ? ( 1'd0 ) : ( n508 ) ;
assign n510 =  ( n166 ) ? ( 1'd0 ) : ( n509 ) ;
assign n511 =  ( n165 ) ? ( 1'd0 ) : ( n510 ) ;
assign n512 =  ( n163 ) ? ( 1'd0 ) : ( n511 ) ;
assign n513 =  ( n158 ) ? ( 1'd0 ) : ( n512 ) ;
assign n514 =  ( n155 ) ? ( 1'd0 ) : ( n513 ) ;
assign n515 =  ( n153 ) ? ( 1'd0 ) : ( n514 ) ;
assign n516 =  ( n133 ) ? ( 1'd0 ) : ( n515 ) ;
assign n517 =  ( n127 ) ? ( 1'd0 ) : ( n516 ) ;
assign n518 =  ( n161 ) ? ( 1'd0 ) : ( n517 ) ;
assign n519 =  ( n160 ) ? ( 1'd0 ) : ( n518 ) ;
assign n520 =  ( n159 ) ? ( 1'd0 ) : ( n519 ) ;
assign n521 =  ( n158 ) ? ( 1'd0 ) : ( n520 ) ;
assign n522 =  ( n157 ) ? ( 1'd0 ) : ( n521 ) ;
assign n523 =  ( n156 ) ? ( 1'd0 ) : ( n522 ) ;
assign n524 =  ( n155 ) ? ( 1'd0 ) : ( n523 ) ;
assign n525 =  ( n154 ) ? ( 1'd0 ) : ( n524 ) ;
assign n526 =  ( n153 ) ? ( 1'd0 ) : ( n525 ) ;
assign n527 =  ( n152 ) ? ( 1'd0 ) : ( n526 ) ;
assign n528 =  ( n151 ) ? ( 1'd0 ) : ( n527 ) ;
assign n529 =  ( n150 ) ? ( 1'd0 ) : ( n528 ) ;
assign n530 =  ( n149 ) ? ( 1'd0 ) : ( n529 ) ;
assign n531 =  ( n148 ) ? ( 1'd0 ) : ( n530 ) ;
assign n532 =  ( n146 ) ? ( 1'd0 ) : ( n531 ) ;
assign n533 =  ( n145 ) ? ( 1'd0 ) : ( n532 ) ;
assign n534 =  ( n144 ) ? ( 1'd0 ) : ( n533 ) ;
assign n535 =  ( n143 ) ? ( 1'd0 ) : ( n534 ) ;
assign n536 =  ( n142 ) ? ( 1'd0 ) : ( n535 ) ;
assign n537 =  ( n141 ) ? ( 1'd0 ) : ( n536 ) ;
assign n538 =  ( n139 ) ? ( 1'd0 ) : ( n537 ) ;
assign n539 =  ( n138 ) ? ( 1'd0 ) : ( n538 ) ;
assign n540 =  ( n137 ) ? ( 1'd0 ) : ( n539 ) ;
assign n541 =  ( n136 ) ? ( 1'd0 ) : ( n540 ) ;
assign n542 =  ( n135 ) ? ( 1'd0 ) : ( n541 ) ;
assign n543 =  ( n134 ) ? ( 1'd0 ) : ( n542 ) ;
assign n544 =  ( n133 ) ? ( 1'd0 ) : ( n543 ) ;
assign n545 =  ( n132 ) ? ( 1'd0 ) : ( n544 ) ;
assign n546 =  ( n131 ) ? ( 1'd0 ) : ( n545 ) ;
assign n547 =  ( n129 ) ? ( 1'd0 ) : ( n546 ) ;
assign n548 =  ( n128 ) ? ( 1'd0 ) : ( n547 ) ;
assign n549 =  ( n127 ) ? ( 1'd0 ) : ( n548 ) ;
assign n550 =  ( n549 ) == ( 1'd1 )  ;
assign n551 =  ( 1'b0 ) | ( n550 )  ;
assign n552 =  ( n115 ) & ( n29 )  ;
assign n553 =  ( n114 ) & ( n4 )  ;
assign n554 =  ( n552 ) | ( n553 )  ;
assign n555 =  ( n116 ) & ( n554 )  ;
assign n556 =  ( n551 ) | ( n555 )  ;
assign n557 =  ( 1'b0 ) ? ( 32'd2048 ) : ( 32'd0 ) ;
assign n558 =  ( 1'b0 ) ? ( 32'd1024 ) : ( n557 ) ;
assign n559 =  ( 1'b0 ) ? ( 32'd512 ) : ( n558 ) ;
assign n560 =  ( 1'b0 ) ? ( 32'd256 ) : ( n559 ) ;
assign n561 =  ( 1'b0 ) ? ( 32'd128 ) : ( n560 ) ;
assign n562 =  ( 1'b0 ) ? ( 32'd64 ) : ( n561 ) ;
assign n563 =  ( 1'b0 ) ? ( 32'd32 ) : ( n562 ) ;
assign n564 =  ( 1'b0 ) ? ( 32'd16 ) : ( n563 ) ;
assign n565 =  ( 1'b0 ) ? ( 32'd8 ) : ( n564 ) ;
assign n566 =  ( n556 ) ? ( 32'd4 ) : ( n565 ) ;
assign n567 =  ( 1'b0 ) ? ( 32'd2 ) : ( n566 ) ;
assign n568__choose_except =  ( n125 ) ? ( 32'd1 ) : ( n567 ) ;
assign n569 = ~ ( medeleg ) ;
assign n570 =  ( n568__choose_except ) & ( n569 )  ;
assign n571 =  ( n570 ) != ( 32'd0 )  ;
assign n572 =  ( n568__choose_except ) & ( medeleg )  ;
assign n573 =  ( n572 ) != ( 32'd0 )  ;
assign n574 =  ( Priv ) > ( 2'd1 )  ;
assign n575 =  ( n573 ) & ( n574 )  ;
assign n576 =  ( n571 ) | ( n575 )  ;
assign n577 =  ( Priv ) <= ( 2'd1 )  ;
assign n578 =  ( n573 ) & ( n577 )  ;
assign n579 = ~ ( n578 ) ;
assign n580 =  ( n576 ) & ( n579 )  ;
assign n581 =  ( n106__take_int_sig ) ? ( n105 ) : ( n580 ) ;
assign n582 =  ( n106__take_int_sig ) ? ( n93 ) : ( n578 ) ;
assign n583 = mstatus[12:11] ;
assign n584 =  ( n583 ) == ( 2'd2 )  ;
assign n585 =  ( n584 ) ? ( 2'd1 ) : ( n583 ) ;
assign n586 = mstatus[8:8] ;
assign n587 =  { ( 1'd0 ) , ( n586 ) }  ;
assign n588 =  ( n115 ) ? ( n585 ) : ( n587 ) ;
assign n589 =  ( n116 ) ? ( n588 ) : ( Priv ) ;
assign n590 =  ( n582 ) ? ( 2'd1 ) : ( n589 ) ;
assign n591 =  ( n581 ) ? ( 2'd3 ) : ( n590 ) ;
assign n592 = ~ ( n106__take_int_sig ) ;
assign n593 = n568__choose_except[0:0] ;
assign n594 = n568__choose_except[1:1] ;
assign n595 =  ( n593 ) | ( n594 )  ;
assign n596 = n568__choose_except[4:4] ;
assign n597 =  ( n595 ) | ( n596 )  ;
assign n598 = n568__choose_except[5:5] ;
assign n599 =  ( n597 ) | ( n598 )  ;
assign n600 = n568__choose_except[6:6] ;
assign n601 =  ( n599 ) | ( n600 )  ;
assign n602 = n568__choose_except[7:7] ;
assign n603 =  ( n601 ) | ( n602 )  ;
assign n604 =  ( n603 ) == ( 1'd1 )  ;
assign n605 =  ( n592 ) & ( n604 )  ;
assign n606 =  ( n605 ) & ( n580 )  ;
assign n607 =  ( n595 ) == ( 1'd1 )  ;
assign n608 =  ( n607 ) ? ( pc ) : ( 32'd0 ) ;
assign n609 =  ( n125 ) | ( 1'b0 )  ;
assign n610 =  ( n609 ) | ( n556 )  ;
assign n611 =  ( n610 ) | ( 1'b0 )  ;
assign n612 =  ( n611 ) | ( 1'b0 )  ;
assign n613 =  ( n612 ) | ( 1'b0 )  ;
assign n614 =  ( n613 ) | ( 1'b0 )  ;
assign n615 =  ( n614 ) | ( 1'b0 )  ;
assign n616 =  ( n615 ) | ( 1'b0 )  ;
assign n617 =  ( n616 ) | ( 1'b0 )  ;
assign n618 =  ( n617 ) | ( 1'b0 )  ;
assign n619 =  ( n618 ) | ( 1'b0 )  ;
assign n620__take_int_or_expt =  ( n619 ) | ( n106__take_int_sig )  ;
assign n621 = ~ ( n620__take_int_or_expt ) ;
assign n622 =  ( n621 ) ? ( mbadaddr ) : ( mbadaddr ) ;
assign n623 =  ( n606 ) ? ( n608 ) : ( n622 ) ;
assign n624 =  ( n581 ) & ( n620__take_int_or_expt )  ;
assign n625 =  ( n97 ) == ( 1'd1 )  ;
assign n626 = n84__int_trap_select[10:10] ;
assign n627 =  ( n626 ) == ( 1'd1 )  ;
assign n628 =  ( n90 ) == ( 1'd1 )  ;
assign n629 = n84__int_trap_select[8:8] ;
assign n630 =  ( n629 ) == ( 1'd1 )  ;
assign n631 =  ( n95 ) == ( 1'd1 )  ;
assign n632 = n84__int_trap_select[6:6] ;
assign n633 =  ( n632 ) == ( 1'd1 )  ;
assign n634 =  ( n87 ) == ( 1'd1 )  ;
assign n635 = n84__int_trap_select[4:4] ;
assign n636 =  ( n635 ) == ( 1'd1 )  ;
assign n637 =  ( n94 ) == ( 1'd1 )  ;
assign n638 = n84__int_trap_select[2:2] ;
assign n639 =  ( n638 ) == ( 1'd1 )  ;
assign n640 =  ( n85 ) == ( 1'd1 )  ;
assign n641 = n84__int_trap_select[0:0] ;
assign n642 =  ( n641 ) == ( 1'd1 )  ;
assign n643 =  ( n642 ) ? ( 32'd0 ) : ( 32'd0 ) ;
assign n644 =  ( n640 ) ? ( 32'd1 ) : ( n643 ) ;
assign n645 =  ( n639 ) ? ( 32'd2 ) : ( n644 ) ;
assign n646 =  ( n637 ) ? ( 32'd3 ) : ( n645 ) ;
assign n647 =  ( n636 ) ? ( 32'd4 ) : ( n646 ) ;
assign n648 =  ( n634 ) ? ( 32'd5 ) : ( n647 ) ;
assign n649 =  ( n633 ) ? ( 32'd6 ) : ( n648 ) ;
assign n650 =  ( n631 ) ? ( 32'd7 ) : ( n649 ) ;
assign n651 =  ( n630 ) ? ( 32'd8 ) : ( n650 ) ;
assign n652 =  ( n628 ) ? ( 32'd9 ) : ( n651 ) ;
assign n653 =  ( n627 ) ? ( 32'd10 ) : ( n652 ) ;
assign n654 =  ( n625 ) ? ( 32'd11 ) : ( n653 ) ;
assign n655 =  ( n654 ) | ( 32'd2147483648 )  ;
assign n656 =  ( 1'b0 ) ? ( 32'd11 ) : ( 32'd12 ) ;
assign n657 =  ( 1'b0 ) ? ( 32'd10 ) : ( n656 ) ;
assign n658 =  ( 1'b0 ) ? ( 32'd9 ) : ( n657 ) ;
assign n659 =  ( 1'b0 ) ? ( 32'd8 ) : ( n658 ) ;
assign n660 =  ( 1'b0 ) ? ( 32'd7 ) : ( n659 ) ;
assign n661 =  ( 1'b0 ) ? ( 32'd6 ) : ( n660 ) ;
assign n662 =  ( 1'b0 ) ? ( 32'd5 ) : ( n661 ) ;
assign n663 =  ( 1'b0 ) ? ( 32'd4 ) : ( n662 ) ;
assign n664 =  ( 1'b0 ) ? ( 32'd3 ) : ( n663 ) ;
assign n665 =  ( n556 ) ? ( 32'd2 ) : ( n664 ) ;
assign n666 =  ( 1'b0 ) ? ( 32'd1 ) : ( n665 ) ;
assign n667__exception_code =  ( n125 ) ? ( 32'd0 ) : ( n666 ) ;
assign n668 =  ( n619 ) ? ( n667__exception_code ) : ( mcause ) ;
assign n669 =  ( n106__take_int_sig ) ? ( n655 ) : ( n668 ) ;
assign n670 =  ( n621 ) ? ( mcause ) : ( mcause ) ;
assign n671 =  ( n624 ) ? ( n669 ) : ( n670 ) ;
assign n672 =  ( n621 ) ? ( medeleg ) : ( medeleg ) ;
assign n673 =  ( pc ) & ( 32'd4294967292 )  ;
assign n674 =  ( n621 ) ? ( mepc ) : ( mepc ) ;
assign n675 =  ( n624 ) ? ( n673 ) : ( n674 ) ;
assign n676 =  ( n621 ) ? ( mideleg ) : ( mideleg ) ;
assign n677 =  ( n621 ) ? ( mie ) : ( mie ) ;
assign n678 =  ( n621 ) ? ( misa ) : ( misa ) ;
assign n679 =  ( n621 ) ? ( mscratch ) : ( mscratch ) ;
assign n680 =  ( n620__take_int_or_expt ) | ( n116 )  ;
assign n681 = ~ ( n582 ) ;
assign n682 =  ( n681 ) & ( n115 )  ;
assign n683 =  ( n682 ) ? ( 2'd0 ) : ( n583 ) ;
assign n684 =  ( n581 ) ? ( Priv ) : ( n683 ) ;
assign n685 = Priv[0:0] ;
assign n686 = ~ ( n581 ) ;
assign n687 =  ( n686 ) & ( n114 )  ;
assign n688 =  ( n687 ) ? ( 1'd0 ) : ( n586 ) ;
assign n689 =  ( n582 ) ? ( n685 ) : ( n688 ) ;
assign n690 =  ( Priv ) == ( 2'd0 )  ;
assign n691 = mstatus[0:0] ;
assign n692 =  ( n690 ) ? ( n691 ) : ( 1'd0 ) ;
assign n693 =  ( n0 ) ? ( n1 ) : ( n692 ) ;
assign n694 =  ( n25 ) ? ( n26 ) : ( n693 ) ;
assign n695 =  ( n681 ) & ( n116 )  ;
assign n696 =  ( n695 ) & ( n115 )  ;
assign n697 = mstatus[7:7] ;
assign n698 =  ( n696 ) ? ( 1'd1 ) : ( n697 ) ;
assign n699 =  ( n581 ) ? ( n694 ) : ( n698 ) ;
assign n700 =  ( n686 ) & ( n116 )  ;
assign n701 =  ( n700 ) & ( n114 )  ;
assign n702 = mstatus[5:5] ;
assign n703 =  ( n701 ) ? ( 1'd1 ) : ( n702 ) ;
assign n704 =  ( n582 ) ? ( n694 ) : ( n703 ) ;
assign n705 =  ( n116 ) & ( n115 )  ;
assign n706 =  ( n583 ) == ( 2'd3 )  ;
assign n707 =  ( n705 ) & ( n706 )  ;
assign n708 =  ( n707 ) ? ( n697 ) : ( n26 ) ;
assign n709 =  ( n582 ) ? ( n26 ) : ( n708 ) ;
assign n710 =  ( n581 ) ? ( 1'd0 ) : ( n709 ) ;
assign n711 =  ( n586 ) == ( 1'd1 )  ;
assign n712 =  ( n114 ) & ( n711 )  ;
assign n713 =  ( n583 ) == ( 2'd1 )  ;
assign n714 =  ( n713 ) | ( n584 )  ;
assign n715 =  ( n115 ) & ( n714 )  ;
assign n716 =  ( n715 ) ? ( n697 ) : ( n1 ) ;
assign n717 =  ( n712 ) ? ( n702 ) : ( n716 ) ;
assign n718 =  ( n116 ) ? ( n717 ) : ( n1 ) ;
assign n719 =  ( n581 ) ? ( n1 ) : ( n718 ) ;
assign n720 =  ( n582 ) ? ( 1'd0 ) : ( n719 ) ;
assign n721 =  { ( n720 ) , ( 1'd0 ) }  ;
assign n722 =  { ( 1'd0 ) , ( n721 ) }  ;
assign n723 =  { ( n710 ) , ( n722 ) }  ;
assign n724 =  { ( 1'd0 ) , ( n723 ) }  ;
assign n725 =  { ( n704 ) , ( n724 ) }  ;
assign n726 =  { ( 1'd0 ) , ( n725 ) }  ;
assign n727 =  { ( n699 ) , ( n726 ) }  ;
assign n728 =  { ( n689 ) , ( n727 ) }  ;
assign n729 =  { ( 2'd0 ) , ( n728 ) }  ;
assign n730 =  { ( n684 ) , ( n729 ) }  ;
assign n731 =  {19'd0 , n730}  ;
assign n732 =  ( n731 ) & ( 32'd6570 )  ;
assign n733 =  ( n621 ) ? ( mstatus ) : ( mstatus ) ;
assign n734 = ~ ( 32'd6570 ) ;
assign n735 =  ( n733 ) & ( n734 )  ;
assign n736 =  ( n732 ) | ( n735 )  ;
assign n737 =  ( n680 ) ? ( n736 ) : ( n733 ) ;
assign n738 =  ( n621 ) ? ( mtvec ) : ( mtvec ) ;
assign n739 =  ( n115 ) ? ( mepc ) : ( sepc ) ;
assign n740 = n113[6:0] ;
assign n741 =  ( n740 ) == ( 7'd103 )  ;
assign n742 = n113[14:12] ;
assign n743 =  ( n742 ) == ( 3'd0 )  ;
assign n744 =  ( n741 ) & ( n743 )  ;
assign n745 = n113[19:15] ;
assign n746 =  ( n745 ) == ( 5'd31 )  ;
assign n747 =  ( n745 ) == ( 5'd30 )  ;
assign n748 =  ( n745 ) == ( 5'd29 )  ;
assign n749 =  ( n745 ) == ( 5'd28 )  ;
assign n750 =  ( n745 ) == ( 5'd27 )  ;
assign n751 =  ( n745 ) == ( 5'd26 )  ;
assign n752 =  ( n745 ) == ( 5'd25 )  ;
assign n753 =  ( n745 ) == ( 5'd24 )  ;
assign n754 =  ( n745 ) == ( 5'd23 )  ;
assign n755 =  ( n745 ) == ( 5'd22 )  ;
assign n756 =  ( n745 ) == ( 5'd21 )  ;
assign n757 =  ( n745 ) == ( 5'd20 )  ;
assign n758 =  ( n745 ) == ( 5'd19 )  ;
assign n759 =  ( n745 ) == ( 5'd18 )  ;
assign n760 =  ( n745 ) == ( 5'd17 )  ;
assign n761 =  ( n745 ) == ( 5'd16 )  ;
assign n762 =  ( n745 ) == ( 5'd15 )  ;
assign n763 =  ( n745 ) == ( 5'd14 )  ;
assign n764 =  ( n745 ) == ( 5'd13 )  ;
assign n765 =  ( n745 ) == ( 5'd12 )  ;
assign n766 =  ( n745 ) == ( 5'd11 )  ;
assign n767 =  ( n745 ) == ( 5'd10 )  ;
assign n768 =  ( n745 ) == ( 5'd9 )  ;
assign n769 =  ( n745 ) == ( 5'd8 )  ;
assign n770 =  ( n745 ) == ( 5'd7 )  ;
assign n771 =  ( n745 ) == ( 5'd6 )  ;
assign n772 =  ( n745 ) == ( 5'd5 )  ;
assign n773 =  ( n745 ) == ( 5'd4 )  ;
assign n774 =  ( n745 ) == ( 5'd3 )  ;
assign n775 =  ( n745 ) == ( 5'd2 )  ;
assign n776 =  ( n745 ) == ( 5'd1 )  ;
assign n777 =  ( n776 ) ? ( x1 ) : ( x0 ) ;
assign n778 =  ( n775 ) ? ( x2 ) : ( n777 ) ;
assign n779 =  ( n774 ) ? ( x3 ) : ( n778 ) ;
assign n780 =  ( n773 ) ? ( x4 ) : ( n779 ) ;
assign n781 =  ( n772 ) ? ( x5 ) : ( n780 ) ;
assign n782 =  ( n771 ) ? ( x6 ) : ( n781 ) ;
assign n783 =  ( n770 ) ? ( x7 ) : ( n782 ) ;
assign n784 =  ( n769 ) ? ( x8 ) : ( n783 ) ;
assign n785 =  ( n768 ) ? ( x9 ) : ( n784 ) ;
assign n786 =  ( n767 ) ? ( x10 ) : ( n785 ) ;
assign n787 =  ( n766 ) ? ( x11 ) : ( n786 ) ;
assign n788 =  ( n765 ) ? ( x12 ) : ( n787 ) ;
assign n789 =  ( n764 ) ? ( x13 ) : ( n788 ) ;
assign n790 =  ( n763 ) ? ( x14 ) : ( n789 ) ;
assign n791 =  ( n762 ) ? ( x15 ) : ( n790 ) ;
assign n792 =  ( n761 ) ? ( x16 ) : ( n791 ) ;
assign n793 =  ( n760 ) ? ( x17 ) : ( n792 ) ;
assign n794 =  ( n759 ) ? ( x18 ) : ( n793 ) ;
assign n795 =  ( n758 ) ? ( x19 ) : ( n794 ) ;
assign n796 =  ( n757 ) ? ( x20 ) : ( n795 ) ;
assign n797 =  ( n756 ) ? ( x21 ) : ( n796 ) ;
assign n798 =  ( n755 ) ? ( x22 ) : ( n797 ) ;
assign n799 =  ( n754 ) ? ( x23 ) : ( n798 ) ;
assign n800 =  ( n753 ) ? ( x24 ) : ( n799 ) ;
assign n801 =  ( n752 ) ? ( x25 ) : ( n800 ) ;
assign n802 =  ( n751 ) ? ( x26 ) : ( n801 ) ;
assign n803 =  ( n750 ) ? ( x27 ) : ( n802 ) ;
assign n804 =  ( n749 ) ? ( x28 ) : ( n803 ) ;
assign n805 =  ( n748 ) ? ( x29 ) : ( n804 ) ;
assign n806 =  ( n747 ) ? ( x30 ) : ( n805 ) ;
assign n807 =  ( n746 ) ? ( x31 ) : ( n806 ) ;
assign n808 = n113[31:20] ;
assign n809 =  { {20{n808[11] }  }, n808}  ;
assign n810 =  ( n807 ) + ( n809 )  ;
assign n811 =  ( n810 ) & ( 32'd4294967294 )  ;
assign n812 =  ( n740 ) == ( 7'd111 )  ;
assign n813 = n113[31:31] ;
assign n814 = n113[19:12] ;
assign n815 = n113[20:20] ;
assign n816 = n113[30:21] ;
assign n817 =  { ( n816 ) , ( 1'd0 ) }  ;
assign n818 =  { ( n815 ) , ( n817 ) }  ;
assign n819 =  { ( n814 ) , ( n818 ) }  ;
assign n820 =  { ( n813 ) , ( n819 ) }  ;
assign n821 =  { {11{n820[20] }  }, n820}  ;
assign n822 =  ( pc ) + ( n821 )  ;
assign n823 =  ( n740 ) == ( 7'd99 )  ;
assign n824 =  ( n742 ) == ( 3'd7 )  ;
assign n825 =  ( n823 ) & ( n824 )  ;
assign n826 = n113[24:20] ;
assign n827 =  ( n826 ) == ( 5'd31 )  ;
assign n828 =  ( n826 ) == ( 5'd30 )  ;
assign n829 =  ( n826 ) == ( 5'd29 )  ;
assign n830 =  ( n826 ) == ( 5'd28 )  ;
assign n831 =  ( n826 ) == ( 5'd27 )  ;
assign n832 =  ( n826 ) == ( 5'd26 )  ;
assign n833 =  ( n826 ) == ( 5'd25 )  ;
assign n834 =  ( n826 ) == ( 5'd24 )  ;
assign n835 =  ( n826 ) == ( 5'd23 )  ;
assign n836 =  ( n826 ) == ( 5'd22 )  ;
assign n837 =  ( n826 ) == ( 5'd21 )  ;
assign n838 =  ( n826 ) == ( 5'd20 )  ;
assign n839 =  ( n826 ) == ( 5'd19 )  ;
assign n840 =  ( n826 ) == ( 5'd18 )  ;
assign n841 =  ( n826 ) == ( 5'd17 )  ;
assign n842 =  ( n826 ) == ( 5'd16 )  ;
assign n843 =  ( n826 ) == ( 5'd15 )  ;
assign n844 =  ( n826 ) == ( 5'd14 )  ;
assign n845 =  ( n826 ) == ( 5'd13 )  ;
assign n846 =  ( n826 ) == ( 5'd12 )  ;
assign n847 =  ( n826 ) == ( 5'd11 )  ;
assign n848 =  ( n826 ) == ( 5'd10 )  ;
assign n849 =  ( n826 ) == ( 5'd9 )  ;
assign n850 =  ( n826 ) == ( 5'd8 )  ;
assign n851 =  ( n826 ) == ( 5'd7 )  ;
assign n852 =  ( n826 ) == ( 5'd6 )  ;
assign n853 =  ( n826 ) == ( 5'd5 )  ;
assign n854 =  ( n826 ) == ( 5'd4 )  ;
assign n855 =  ( n826 ) == ( 5'd3 )  ;
assign n856 =  ( n826 ) == ( 5'd2 )  ;
assign n857 =  ( n826 ) == ( 5'd1 )  ;
assign n858 =  ( n857 ) ? ( x1 ) : ( x0 ) ;
assign n859 =  ( n856 ) ? ( x2 ) : ( n858 ) ;
assign n860 =  ( n855 ) ? ( x3 ) : ( n859 ) ;
assign n861 =  ( n854 ) ? ( x4 ) : ( n860 ) ;
assign n862 =  ( n853 ) ? ( x5 ) : ( n861 ) ;
assign n863 =  ( n852 ) ? ( x6 ) : ( n862 ) ;
assign n864 =  ( n851 ) ? ( x7 ) : ( n863 ) ;
assign n865 =  ( n850 ) ? ( x8 ) : ( n864 ) ;
assign n866 =  ( n849 ) ? ( x9 ) : ( n865 ) ;
assign n867 =  ( n848 ) ? ( x10 ) : ( n866 ) ;
assign n868 =  ( n847 ) ? ( x11 ) : ( n867 ) ;
assign n869 =  ( n846 ) ? ( x12 ) : ( n868 ) ;
assign n870 =  ( n845 ) ? ( x13 ) : ( n869 ) ;
assign n871 =  ( n844 ) ? ( x14 ) : ( n870 ) ;
assign n872 =  ( n843 ) ? ( x15 ) : ( n871 ) ;
assign n873 =  ( n842 ) ? ( x16 ) : ( n872 ) ;
assign n874 =  ( n841 ) ? ( x17 ) : ( n873 ) ;
assign n875 =  ( n840 ) ? ( x18 ) : ( n874 ) ;
assign n876 =  ( n839 ) ? ( x19 ) : ( n875 ) ;
assign n877 =  ( n838 ) ? ( x20 ) : ( n876 ) ;
assign n878 =  ( n837 ) ? ( x21 ) : ( n877 ) ;
assign n879 =  ( n836 ) ? ( x22 ) : ( n878 ) ;
assign n880 =  ( n835 ) ? ( x23 ) : ( n879 ) ;
assign n881 =  ( n834 ) ? ( x24 ) : ( n880 ) ;
assign n882 =  ( n833 ) ? ( x25 ) : ( n881 ) ;
assign n883 =  ( n832 ) ? ( x26 ) : ( n882 ) ;
assign n884 =  ( n831 ) ? ( x27 ) : ( n883 ) ;
assign n885 =  ( n830 ) ? ( x28 ) : ( n884 ) ;
assign n886 =  ( n829 ) ? ( x29 ) : ( n885 ) ;
assign n887 =  ( n828 ) ? ( x30 ) : ( n886 ) ;
assign n888 =  ( n827 ) ? ( x31 ) : ( n887 ) ;
assign n889 =  ( n807 ) >= ( n888 )  ;
assign n890 = n113[7:7] ;
assign n891 = n113[30:25] ;
assign n892 = n113[11:8] ;
assign n893 =  { ( n892 ) , ( 1'd0 ) }  ;
assign n894 =  { ( n891 ) , ( n893 ) }  ;
assign n895 =  { ( n890 ) , ( n894 ) }  ;
assign n896 =  { ( n813 ) , ( n895 ) }  ;
assign n897 =  { {19{n896[12] }  }, n896}  ;
assign n898 =  ( pc ) + ( n897 )  ;
assign n899 =  ( pc ) + ( 32'd4 )  ;
assign n900 =  ( n889 ) ? ( n898 ) : ( n899 ) ;
assign n901 =  ( n742 ) == ( 3'd5 )  ;
assign n902 =  ( n823 ) & ( n901 )  ;
assign n903 =  $signed( n807 ) >= $signed( n888 )  ;
assign n904 =  ( n903 ) ? ( n898 ) : ( n899 ) ;
assign n905 =  ( n742 ) == ( 3'd6 )  ;
assign n906 =  ( n823 ) & ( n905 )  ;
assign n907 =  ( n807 ) < ( n888 )  ;
assign n908 =  ( n907 ) ? ( n898 ) : ( n899 ) ;
assign n909 =  ( n742 ) == ( 3'd4 )  ;
assign n910 =  ( n823 ) & ( n909 )  ;
assign n911 =  $signed( n807 ) < $signed( n888 )  ;
assign n912 =  ( n911 ) ? ( n898 ) : ( n899 ) ;
assign n913 =  ( n742 ) == ( 3'd1 )  ;
assign n914 =  ( n823 ) & ( n913 )  ;
assign n915 =  ( n807 ) != ( n888 )  ;
assign n916 =  ( n915 ) ? ( n898 ) : ( n899 ) ;
assign n917 =  ( n823 ) & ( n743 )  ;
assign n918 =  ( n807 ) == ( n888 )  ;
assign n919 =  ( n918 ) ? ( n898 ) : ( n899 ) ;
assign n920 =  ( n740 ) == ( 7'd51 )  ;
assign n921 =  ( n920 ) & ( n901 )  ;
assign n922 = n113[31:25] ;
assign n923 =  ( n922 ) == ( 7'd32 )  ;
assign n924 =  ( n921 ) & ( n923 )  ;
assign n925 =  ( n920 ) & ( n743 )  ;
assign n926 =  ( n925 ) & ( n923 )  ;
assign n927 =  ( n922 ) == ( 7'd0 )  ;
assign n928 =  ( n921 ) & ( n927 )  ;
assign n929 =  ( n920 ) & ( n913 )  ;
assign n930 =  ( n929 ) & ( n927 )  ;
assign n931 =  ( n920 ) & ( n909 )  ;
assign n932 =  ( n931 ) & ( n927 )  ;
assign n933 =  ( n920 ) & ( n905 )  ;
assign n934 =  ( n933 ) & ( n927 )  ;
assign n935 =  ( n920 ) & ( n824 )  ;
assign n936 =  ( n935 ) & ( n927 )  ;
assign n937 =  ( n742 ) == ( 3'd3 )  ;
assign n938 =  ( n920 ) & ( n937 )  ;
assign n939 =  ( n938 ) & ( n927 )  ;
assign n940 =  ( n742 ) == ( 3'd2 )  ;
assign n941 =  ( n920 ) & ( n940 )  ;
assign n942 =  ( n941 ) & ( n927 )  ;
assign n943 =  ( n925 ) & ( n927 )  ;
assign n944 =  ( n740 ) == ( 7'd19 )  ;
assign n945 =  ( n944 ) & ( n901 )  ;
assign n946 =  ( n945 ) & ( n923 )  ;
assign n947 =  ( n945 ) & ( n927 )  ;
assign n948 =  ( n944 ) & ( n913 )  ;
assign n949 =  ( n948 ) & ( n927 )  ;
assign n950 =  ( n944 ) & ( n909 )  ;
assign n951 =  ( n944 ) & ( n905 )  ;
assign n952 =  ( n944 ) & ( n824 )  ;
assign n953 =  ( n944 ) & ( n937 )  ;
assign n954 =  ( n944 ) & ( n940 )  ;
assign n955 =  ( n944 ) & ( n743 )  ;
assign n956 =  ( n740 ) == ( 7'd23 )  ;
assign n957 =  ( n740 ) == ( 7'd55 )  ;
assign n958 =  ( n740 ) == ( 7'd35 )  ;
assign n959 =  ( n958 ) & ( n940 )  ;
assign n960 =  ( n958 ) & ( n913 )  ;
assign n961 =  ( n958 ) & ( n743 )  ;
assign n962 =  ( n740 ) == ( 7'd3 )  ;
assign n963 =  ( n962 ) & ( n901 )  ;
assign n964 =  ( n962 ) & ( n909 )  ;
assign n965 =  ( n962 ) & ( n743 )  ;
assign n966 =  ( n962 ) & ( n913 )  ;
assign n967 =  ( n962 ) & ( n940 )  ;
assign n968 =  ( n966 ) | ( n967 )  ;
assign n969 =  ( n965 ) | ( n968 )  ;
assign n970 =  ( n964 ) | ( n969 )  ;
assign n971 =  ( n963 ) | ( n970 )  ;
assign n972 =  ( n961 ) | ( n971 )  ;
assign n973 =  ( n960 ) | ( n972 )  ;
assign n974 =  ( n959 ) | ( n973 )  ;
assign n975 =  ( n957 ) | ( n974 )  ;
assign n976 =  ( n956 ) | ( n975 )  ;
assign n977 =  ( n955 ) | ( n976 )  ;
assign n978 =  ( n954 ) | ( n977 )  ;
assign n979 =  ( n953 ) | ( n978 )  ;
assign n980 =  ( n952 ) | ( n979 )  ;
assign n981 =  ( n951 ) | ( n980 )  ;
assign n982 =  ( n950 ) | ( n981 )  ;
assign n983 =  ( n949 ) | ( n982 )  ;
assign n984 =  ( n947 ) | ( n983 )  ;
assign n985 =  ( n946 ) | ( n984 )  ;
assign n986 =  ( n943 ) | ( n985 )  ;
assign n987 =  ( n942 ) | ( n986 )  ;
assign n988 =  ( n939 ) | ( n987 )  ;
assign n989 =  ( n936 ) | ( n988 )  ;
assign n990 =  ( n934 ) | ( n989 )  ;
assign n991 =  ( n932 ) | ( n990 )  ;
assign n992 =  ( n930 ) | ( n991 )  ;
assign n993 =  ( n928 ) | ( n992 )  ;
assign n994 =  ( n926 ) | ( n993 )  ;
assign n995 =  ( n924 ) | ( n994 )  ;
assign n996 =  ( n995 ) ? ( n899 ) : ( pc ) ;
assign n997 =  ( n917 ) ? ( n919 ) : ( n996 ) ;
assign n998 =  ( n914 ) ? ( n916 ) : ( n997 ) ;
assign n999 =  ( n910 ) ? ( n912 ) : ( n998 ) ;
assign n1000 =  ( n906 ) ? ( n908 ) : ( n999 ) ;
assign n1001 =  ( n902 ) ? ( n904 ) : ( n1000 ) ;
assign n1002 =  ( n825 ) ? ( n900 ) : ( n1001 ) ;
assign n1003 =  ( n812 ) ? ( n822 ) : ( n1002 ) ;
assign n1004 =  ( n744 ) ? ( n811 ) : ( n1003 ) ;
assign n1005 =  ( n116 ) ? ( n739 ) : ( n1004 ) ;
assign n1006 =  ( n582 ) ? ( stvec ) : ( n1005 ) ;
assign n1007 =  ( n581 ) ? ( mtvec ) : ( n1006 ) ;
assign n1008 =  ( n605 ) & ( n578 )  ;
assign n1009 =  ( n621 ) ? ( sbadaddr ) : ( sbadaddr ) ;
assign n1010 =  ( n1008 ) ? ( n608 ) : ( n1009 ) ;
assign n1011 =  ( n582 ) & ( n620__take_int_or_expt )  ;
assign n1012 =  ( n619 ) ? ( n667__exception_code ) : ( scause ) ;
assign n1013 =  ( n106__take_int_sig ) ? ( n655 ) : ( n1012 ) ;
assign n1014 =  ( n621 ) ? ( scause ) : ( scause ) ;
assign n1015 =  ( n1011 ) ? ( n1013 ) : ( n1014 ) ;
assign n1016 =  ( n621 ) ? ( sepc ) : ( sepc ) ;
assign n1017 =  ( n1011 ) ? ( n673 ) : ( n1016 ) ;
assign n1018 =  ( n621 ) ? ( sptbr ) : ( sptbr ) ;
assign n1019 =  ( n621 ) ? ( sscratch ) : ( sscratch ) ;
assign n1020 =  ( n621 ) ? ( stvec ) : ( stvec ) ;
assign n1021 = n113[11:7] ;
assign n1022 =  ( n1021 ) == ( 5'd1 )  ;
assign n1023 = n888[4:0] ;
assign n1024 =  {27'd0 , n1023}  ;
assign n1025 =  ( $signed( n807 ) >>> ( n1024 ))  ;
assign n1026 =  ( n1022 ) ? ( n1025 ) : ( x1 ) ;
assign n1027 =  ( n807 ) - ( n888 )  ;
assign n1028 =  ( n1022 ) ? ( n1027 ) : ( x1 ) ;
assign n1029 =  ( ( n807 ) >> ( n1024 ))  ;
assign n1030 =  ( n1022 ) ? ( n1029 ) : ( x1 ) ;
assign n1031 =  ( n807 ) << ( n1024 )  ;
assign n1032 =  ( n1022 ) ? ( n1031 ) : ( x1 ) ;
assign n1033 =  ( n807 ) ^ ( n888 )  ;
assign n1034 =  ( n1022 ) ? ( n1033 ) : ( x1 ) ;
assign n1035 =  ( n807 ) | ( n888 )  ;
assign n1036 =  ( n1022 ) ? ( n1035 ) : ( x1 ) ;
assign n1037 =  ( n807 ) & ( n888 )  ;
assign n1038 =  ( n1022 ) ? ( n1037 ) : ( x1 ) ;
assign n1039 =  ( n907 ) ? ( 32'd1 ) : ( 32'd0 ) ;
assign n1040 =  ( n1022 ) ? ( n1039 ) : ( x1 ) ;
assign n1041 =  ( n911 ) ? ( 32'd1 ) : ( 32'd0 ) ;
assign n1042 =  ( n1022 ) ? ( n1041 ) : ( x1 ) ;
assign n1043 =  ( n807 ) + ( n888 )  ;
assign n1044 =  ( n1022 ) ? ( n1043 ) : ( x1 ) ;
assign n1045 =  {27'd0 , n826}  ;
assign n1046 =  ( $signed( n807 ) >>> ( n1045 ))  ;
assign n1047 =  ( n1022 ) ? ( n1046 ) : ( x1 ) ;
assign n1048 =  ( ( n807 ) >> ( n1045 ))  ;
assign n1049 =  ( n1022 ) ? ( n1048 ) : ( x1 ) ;
assign n1050 =  ( n807 ) << ( n1045 )  ;
assign n1051 =  ( n1022 ) ? ( n1050 ) : ( x1 ) ;
assign n1052 = n809 ;
assign n1053 =  ( n807 ) ^ ( n1052 )  ;
assign n1054 =  ( n1022 ) ? ( n1053 ) : ( x1 ) ;
assign n1055 = n809 ;
assign n1056 =  ( n807 ) | ( n1055 )  ;
assign n1057 =  ( n1022 ) ? ( n1056 ) : ( x1 ) ;
assign n1058 =  ( n807 ) & ( n1052 )  ;
assign n1059 =  ( n1022 ) ? ( n1058 ) : ( x1 ) ;
assign n1060 =  ( n807 ) < ( n1055 )  ;
assign n1061 =  ( n1060 ) ? ( 32'd1 ) : ( 32'd0 ) ;
assign n1062 =  ( n1022 ) ? ( n1061 ) : ( x1 ) ;
assign n1063 =  $signed( n807 ) < $signed( n1052 )  ;
assign n1064 =  ( n1063 ) ? ( 32'd1 ) : ( 32'd0 ) ;
assign n1065 =  ( n1022 ) ? ( n1064 ) : ( x1 ) ;
assign n1066 =  ( n807 ) + ( n1052 )  ;
assign n1067 =  ( n1022 ) ? ( n1066 ) : ( x1 ) ;
assign n1068 =  ( n744 ) | ( n812 )  ;
assign n1069 =  ( n1022 ) ? ( n899 ) : ( x1 ) ;
assign n1070 = n113[31:12] ;
assign n1071 =  { ( n1070 ) , ( 12'd0 ) }  ;
assign n1072 =  ( n1071 ) + ( pc )  ;
assign n1073 =  ( n1022 ) ? ( n1072 ) : ( x1 ) ;
assign n1074 =  ( n1022 ) ? ( n1071 ) : ( x1 ) ;
assign n1075 = n810[1:0] ;
assign n1076 =  ( n1075 ) == ( 2'd0 )  ;
assign n1077 = n810[31:2] ;
assign n1078 =  {2'd0 , n1077}  ;
assign mem_addr_n1079 = n1078 ;
assign n1081 = mem_data_n1080 ;
assign n1082 = n1081[15:0] ;
assign n1083 =  {16'd0 , n1082}  ;
assign n1084 =  ( n1075 ) == ( 2'd1 )  ;
assign n1085 = n1081[15:8] ;
assign n1086 =  {24'd0 , n1085}  ;
assign n1087 =  ( n1075 ) == ( 2'd2 )  ;
assign n1088 = n1081[31:16] ;
assign n1089 =  {16'd0 , n1088}  ;
assign n1090 =  ( n1075 ) == ( 2'd3 )  ;
assign n1091 = n1081[31:24] ;
assign n1092 =  {24'd0 , n1091}  ;
assign n1093 = n1081[31:0] ;
assign n1094 =  ( n1090 ) ? ( n1092 ) : ( n1093 ) ;
assign n1095 =  ( n1087 ) ? ( n1089 ) : ( n1094 ) ;
assign n1096 =  ( n1084 ) ? ( n1086 ) : ( n1095 ) ;
assign n1097 =  ( n1076 ) ? ( n1083 ) : ( n1096 ) ;
assign n1098 =  ( n1022 ) ? ( n1097 ) : ( x1 ) ;
assign n1099 = n1081[7:0] ;
assign n1100 =  {24'd0 , n1099}  ;
assign n1101 = n1081[23:16] ;
assign n1102 =  {24'd0 , n1101}  ;
assign n1103 =  ( n1087 ) ? ( n1102 ) : ( n1094 ) ;
assign n1104 =  ( n1084 ) ? ( n1086 ) : ( n1103 ) ;
assign n1105 =  ( n1076 ) ? ( n1100 ) : ( n1104 ) ;
assign n1106 =  ( n1022 ) ? ( n1105 ) : ( x1 ) ;
assign n1107 =  { {24{n1099[7] }  }, n1099}  ;
assign n1108 =  { {24{n1085[7] }  }, n1085}  ;
assign n1109 =  { {24{n1101[7] }  }, n1101}  ;
assign n1110 =  { {24{n1091[7] }  }, n1091}  ;
assign n1111 =  ( n1090 ) ? ( n1110 ) : ( n1093 ) ;
assign n1112 =  ( n1087 ) ? ( n1109 ) : ( n1111 ) ;
assign n1113 =  ( n1084 ) ? ( n1108 ) : ( n1112 ) ;
assign n1114 =  ( n1076 ) ? ( n1107 ) : ( n1113 ) ;
assign n1115 =  ( n1022 ) ? ( n1114 ) : ( x1 ) ;
assign n1116 =  { {16{n1082[15] }  }, n1082}  ;
assign n1117 =  { {16{n1088[15] }  }, n1088}  ;
assign n1118 =  ( n1087 ) ? ( n1117 ) : ( n1094 ) ;
assign n1119 =  ( n1084 ) ? ( n1086 ) : ( n1118 ) ;
assign n1120 =  ( n1076 ) ? ( n1116 ) : ( n1119 ) ;
assign n1121 =  ( n1022 ) ? ( n1120 ) : ( x1 ) ;
assign n1122 =  ( n1076 ) ? ( n1093 ) : ( n1104 ) ;
assign n1123 =  ( n1022 ) ? ( n1122 ) : ( x1 ) ;
assign n1124 =  ( n967 ) ? ( n1123 ) : ( x1 ) ;
assign n1125 =  ( n966 ) ? ( n1121 ) : ( n1124 ) ;
assign n1126 =  ( n965 ) ? ( n1115 ) : ( n1125 ) ;
assign n1127 =  ( n964 ) ? ( n1106 ) : ( n1126 ) ;
assign n1128 =  ( n963 ) ? ( n1098 ) : ( n1127 ) ;
assign n1129 =  ( n957 ) ? ( n1074 ) : ( n1128 ) ;
assign n1130 =  ( n956 ) ? ( n1073 ) : ( n1129 ) ;
assign n1131 =  ( n1068 ) ? ( n1069 ) : ( n1130 ) ;
assign n1132 =  ( n955 ) ? ( n1067 ) : ( n1131 ) ;
assign n1133 =  ( n954 ) ? ( n1065 ) : ( n1132 ) ;
assign n1134 =  ( n953 ) ? ( n1062 ) : ( n1133 ) ;
assign n1135 =  ( n952 ) ? ( n1059 ) : ( n1134 ) ;
assign n1136 =  ( n951 ) ? ( n1057 ) : ( n1135 ) ;
assign n1137 =  ( n950 ) ? ( n1054 ) : ( n1136 ) ;
assign n1138 =  ( n949 ) ? ( n1051 ) : ( n1137 ) ;
assign n1139 =  ( n947 ) ? ( n1049 ) : ( n1138 ) ;
assign n1140 =  ( n946 ) ? ( n1047 ) : ( n1139 ) ;
assign n1141 =  ( n943 ) ? ( n1044 ) : ( n1140 ) ;
assign n1142 =  ( n942 ) ? ( n1042 ) : ( n1141 ) ;
assign n1143 =  ( n939 ) ? ( n1040 ) : ( n1142 ) ;
assign n1144 =  ( n936 ) ? ( n1038 ) : ( n1143 ) ;
assign n1145 =  ( n934 ) ? ( n1036 ) : ( n1144 ) ;
assign n1146 =  ( n932 ) ? ( n1034 ) : ( n1145 ) ;
assign n1147 =  ( n930 ) ? ( n1032 ) : ( n1146 ) ;
assign n1148 =  ( n928 ) ? ( n1030 ) : ( n1147 ) ;
assign n1149 =  ( n926 ) ? ( n1028 ) : ( n1148 ) ;
assign n1150 =  ( n924 ) ? ( n1026 ) : ( n1149 ) ;
assign n1151 =  ( n621 ) ? ( n1150 ) : ( x1 ) ;
assign n1152 =  ( n1021 ) == ( 5'd10 )  ;
assign n1153 =  ( n1152 ) ? ( n1025 ) : ( x10 ) ;
assign n1154 =  ( n1152 ) ? ( n1027 ) : ( x10 ) ;
assign n1155 =  ( n1152 ) ? ( n1029 ) : ( x10 ) ;
assign n1156 =  ( n1152 ) ? ( n1031 ) : ( x10 ) ;
assign n1157 =  ( n1152 ) ? ( n1033 ) : ( x10 ) ;
assign n1158 =  ( n1152 ) ? ( n1035 ) : ( x10 ) ;
assign n1159 =  ( n1152 ) ? ( n1037 ) : ( x10 ) ;
assign n1160 =  ( n1152 ) ? ( n1039 ) : ( x10 ) ;
assign n1161 =  ( n1152 ) ? ( n1041 ) : ( x10 ) ;
assign n1162 =  ( n1152 ) ? ( n1043 ) : ( x10 ) ;
assign n1163 =  ( n1152 ) ? ( n1046 ) : ( x10 ) ;
assign n1164 =  ( n1152 ) ? ( n1048 ) : ( x10 ) ;
assign n1165 =  ( n1152 ) ? ( n1050 ) : ( x10 ) ;
assign n1166 =  ( n1152 ) ? ( n1053 ) : ( x10 ) ;
assign n1167 =  ( n807 ) | ( n1052 )  ;
assign n1168 =  ( n1152 ) ? ( n1167 ) : ( x10 ) ;
assign n1169 =  ( n1152 ) ? ( n1058 ) : ( x10 ) ;
assign n1170 =  ( n1152 ) ? ( n1061 ) : ( x10 ) ;
assign n1171 =  ( n1152 ) ? ( n1064 ) : ( x10 ) ;
assign n1172 =  ( n1152 ) ? ( n1066 ) : ( x10 ) ;
assign n1173 =  ( n1152 ) ? ( n899 ) : ( x10 ) ;
assign n1174 =  ( n1152 ) ? ( n1072 ) : ( x10 ) ;
assign n1175 =  ( n1152 ) ? ( n1071 ) : ( x10 ) ;
assign n1176 =  ( n1152 ) ? ( n1097 ) : ( x10 ) ;
assign n1177 =  ( n1152 ) ? ( n1105 ) : ( x10 ) ;
assign n1178 =  ( n1152 ) ? ( n1114 ) : ( x10 ) ;
assign n1179 =  ( n1152 ) ? ( n1120 ) : ( x10 ) ;
assign n1180 =  ( n1152 ) ? ( n1122 ) : ( x10 ) ;
assign n1181 =  ( n967 ) ? ( n1180 ) : ( x10 ) ;
assign n1182 =  ( n966 ) ? ( n1179 ) : ( n1181 ) ;
assign n1183 =  ( n965 ) ? ( n1178 ) : ( n1182 ) ;
assign n1184 =  ( n964 ) ? ( n1177 ) : ( n1183 ) ;
assign n1185 =  ( n963 ) ? ( n1176 ) : ( n1184 ) ;
assign n1186 =  ( n957 ) ? ( n1175 ) : ( n1185 ) ;
assign n1187 =  ( n956 ) ? ( n1174 ) : ( n1186 ) ;
assign n1188 =  ( n1068 ) ? ( n1173 ) : ( n1187 ) ;
assign n1189 =  ( n955 ) ? ( n1172 ) : ( n1188 ) ;
assign n1190 =  ( n954 ) ? ( n1171 ) : ( n1189 ) ;
assign n1191 =  ( n953 ) ? ( n1170 ) : ( n1190 ) ;
assign n1192 =  ( n952 ) ? ( n1169 ) : ( n1191 ) ;
assign n1193 =  ( n951 ) ? ( n1168 ) : ( n1192 ) ;
assign n1194 =  ( n950 ) ? ( n1166 ) : ( n1193 ) ;
assign n1195 =  ( n949 ) ? ( n1165 ) : ( n1194 ) ;
assign n1196 =  ( n947 ) ? ( n1164 ) : ( n1195 ) ;
assign n1197 =  ( n946 ) ? ( n1163 ) : ( n1196 ) ;
assign n1198 =  ( n943 ) ? ( n1162 ) : ( n1197 ) ;
assign n1199 =  ( n942 ) ? ( n1161 ) : ( n1198 ) ;
assign n1200 =  ( n939 ) ? ( n1160 ) : ( n1199 ) ;
assign n1201 =  ( n936 ) ? ( n1159 ) : ( n1200 ) ;
assign n1202 =  ( n934 ) ? ( n1158 ) : ( n1201 ) ;
assign n1203 =  ( n932 ) ? ( n1157 ) : ( n1202 ) ;
assign n1204 =  ( n930 ) ? ( n1156 ) : ( n1203 ) ;
assign n1205 =  ( n928 ) ? ( n1155 ) : ( n1204 ) ;
assign n1206 =  ( n926 ) ? ( n1154 ) : ( n1205 ) ;
assign n1207 =  ( n924 ) ? ( n1153 ) : ( n1206 ) ;
assign n1208 =  ( n621 ) ? ( n1207 ) : ( x10 ) ;
assign n1209 =  ( n1021 ) == ( 5'd11 )  ;
assign n1210 =  ( n1209 ) ? ( n1025 ) : ( x11 ) ;
assign n1211 =  ( n1209 ) ? ( n1027 ) : ( x11 ) ;
assign n1212 =  ( n1209 ) ? ( n1029 ) : ( x11 ) ;
assign n1213 =  ( n1209 ) ? ( n1031 ) : ( x11 ) ;
assign n1214 =  ( n1209 ) ? ( n1033 ) : ( x11 ) ;
assign n1215 =  ( n1209 ) ? ( n1035 ) : ( x11 ) ;
assign n1216 =  ( n1209 ) ? ( n1037 ) : ( x11 ) ;
assign n1217 =  ( n1209 ) ? ( n1039 ) : ( x11 ) ;
assign n1218 =  ( n1209 ) ? ( n1041 ) : ( x11 ) ;
assign n1219 =  ( n1209 ) ? ( n1043 ) : ( x11 ) ;
assign n1220 =  ( n1209 ) ? ( n1046 ) : ( x11 ) ;
assign n1221 =  ( n1209 ) ? ( n1048 ) : ( x11 ) ;
assign n1222 =  ( n1209 ) ? ( n1050 ) : ( x11 ) ;
assign n1223 =  ( n1209 ) ? ( n1053 ) : ( x11 ) ;
assign n1224 =  ( n1209 ) ? ( n1167 ) : ( x11 ) ;
assign n1225 =  ( n1209 ) ? ( n1058 ) : ( x11 ) ;
assign n1226 =  ( n1209 ) ? ( n1061 ) : ( x11 ) ;
assign n1227 =  ( n1209 ) ? ( n1064 ) : ( x11 ) ;
assign n1228 =  ( n1209 ) ? ( n1066 ) : ( x11 ) ;
assign n1229 =  ( n1209 ) ? ( n899 ) : ( x11 ) ;
assign n1230 =  ( n1209 ) ? ( n1072 ) : ( x11 ) ;
assign n1231 =  ( n1209 ) ? ( n1071 ) : ( x11 ) ;
assign n1232 =  ( n1209 ) ? ( n1097 ) : ( x11 ) ;
assign n1233 =  ( n1209 ) ? ( n1105 ) : ( x11 ) ;
assign n1234 =  ( n1209 ) ? ( n1114 ) : ( x11 ) ;
assign n1235 =  ( n1209 ) ? ( n1120 ) : ( x11 ) ;
assign n1236 =  ( n1209 ) ? ( n1122 ) : ( x11 ) ;
assign n1237 =  ( n967 ) ? ( n1236 ) : ( x11 ) ;
assign n1238 =  ( n966 ) ? ( n1235 ) : ( n1237 ) ;
assign n1239 =  ( n965 ) ? ( n1234 ) : ( n1238 ) ;
assign n1240 =  ( n964 ) ? ( n1233 ) : ( n1239 ) ;
assign n1241 =  ( n963 ) ? ( n1232 ) : ( n1240 ) ;
assign n1242 =  ( n957 ) ? ( n1231 ) : ( n1241 ) ;
assign n1243 =  ( n956 ) ? ( n1230 ) : ( n1242 ) ;
assign n1244 =  ( n1068 ) ? ( n1229 ) : ( n1243 ) ;
assign n1245 =  ( n955 ) ? ( n1228 ) : ( n1244 ) ;
assign n1246 =  ( n954 ) ? ( n1227 ) : ( n1245 ) ;
assign n1247 =  ( n953 ) ? ( n1226 ) : ( n1246 ) ;
assign n1248 =  ( n952 ) ? ( n1225 ) : ( n1247 ) ;
assign n1249 =  ( n951 ) ? ( n1224 ) : ( n1248 ) ;
assign n1250 =  ( n950 ) ? ( n1223 ) : ( n1249 ) ;
assign n1251 =  ( n949 ) ? ( n1222 ) : ( n1250 ) ;
assign n1252 =  ( n947 ) ? ( n1221 ) : ( n1251 ) ;
assign n1253 =  ( n946 ) ? ( n1220 ) : ( n1252 ) ;
assign n1254 =  ( n943 ) ? ( n1219 ) : ( n1253 ) ;
assign n1255 =  ( n942 ) ? ( n1218 ) : ( n1254 ) ;
assign n1256 =  ( n939 ) ? ( n1217 ) : ( n1255 ) ;
assign n1257 =  ( n936 ) ? ( n1216 ) : ( n1256 ) ;
assign n1258 =  ( n934 ) ? ( n1215 ) : ( n1257 ) ;
assign n1259 =  ( n932 ) ? ( n1214 ) : ( n1258 ) ;
assign n1260 =  ( n930 ) ? ( n1213 ) : ( n1259 ) ;
assign n1261 =  ( n928 ) ? ( n1212 ) : ( n1260 ) ;
assign n1262 =  ( n926 ) ? ( n1211 ) : ( n1261 ) ;
assign n1263 =  ( n924 ) ? ( n1210 ) : ( n1262 ) ;
assign n1264 =  ( n621 ) ? ( n1263 ) : ( x11 ) ;
assign n1265 =  ( n1021 ) == ( 5'd12 )  ;
assign n1266 =  ( n1265 ) ? ( n1025 ) : ( x12 ) ;
assign n1267 =  ( n1265 ) ? ( n1027 ) : ( x12 ) ;
assign n1268 =  ( n1265 ) ? ( n1029 ) : ( x12 ) ;
assign n1269 =  ( n1265 ) ? ( n1031 ) : ( x12 ) ;
assign n1270 =  ( n1265 ) ? ( n1033 ) : ( x12 ) ;
assign n1271 =  ( n1265 ) ? ( n1035 ) : ( x12 ) ;
assign n1272 =  ( n1265 ) ? ( n1037 ) : ( x12 ) ;
assign n1273 =  ( n1265 ) ? ( n1039 ) : ( x12 ) ;
assign n1274 =  ( n1265 ) ? ( n1041 ) : ( x12 ) ;
assign n1275 =  ( n1265 ) ? ( n1043 ) : ( x12 ) ;
assign n1276 =  ( n1265 ) ? ( n1046 ) : ( x12 ) ;
assign n1277 =  ( n1265 ) ? ( n1048 ) : ( x12 ) ;
assign n1278 =  ( n1265 ) ? ( n1050 ) : ( x12 ) ;
assign n1279 =  ( n1265 ) ? ( n1053 ) : ( x12 ) ;
assign n1280 =  ( n1265 ) ? ( n1167 ) : ( x12 ) ;
assign n1281 =  ( n1265 ) ? ( n1058 ) : ( x12 ) ;
assign n1282 =  ( n807 ) < ( n1052 )  ;
assign n1283 =  ( n1282 ) ? ( 32'd1 ) : ( 32'd0 ) ;
assign n1284 =  ( n1265 ) ? ( n1283 ) : ( x12 ) ;
assign n1285 =  ( n1265 ) ? ( n1064 ) : ( x12 ) ;
assign n1286 =  ( n1265 ) ? ( n1066 ) : ( x12 ) ;
assign n1287 =  ( n1265 ) ? ( n899 ) : ( x12 ) ;
assign n1288 =  ( n1265 ) ? ( n1072 ) : ( x12 ) ;
assign n1289 =  ( n1265 ) ? ( n1071 ) : ( x12 ) ;
assign n1290 =  ( n1265 ) ? ( n1097 ) : ( x12 ) ;
assign n1291 =  ( n1265 ) ? ( n1105 ) : ( x12 ) ;
assign n1292 =  ( n1265 ) ? ( n1114 ) : ( x12 ) ;
assign n1293 =  ( n1265 ) ? ( n1120 ) : ( x12 ) ;
assign n1294 =  ( n1265 ) ? ( n1122 ) : ( x12 ) ;
assign n1295 =  ( n967 ) ? ( n1294 ) : ( x12 ) ;
assign n1296 =  ( n966 ) ? ( n1293 ) : ( n1295 ) ;
assign n1297 =  ( n965 ) ? ( n1292 ) : ( n1296 ) ;
assign n1298 =  ( n964 ) ? ( n1291 ) : ( n1297 ) ;
assign n1299 =  ( n963 ) ? ( n1290 ) : ( n1298 ) ;
assign n1300 =  ( n957 ) ? ( n1289 ) : ( n1299 ) ;
assign n1301 =  ( n956 ) ? ( n1288 ) : ( n1300 ) ;
assign n1302 =  ( n1068 ) ? ( n1287 ) : ( n1301 ) ;
assign n1303 =  ( n955 ) ? ( n1286 ) : ( n1302 ) ;
assign n1304 =  ( n954 ) ? ( n1285 ) : ( n1303 ) ;
assign n1305 =  ( n953 ) ? ( n1284 ) : ( n1304 ) ;
assign n1306 =  ( n952 ) ? ( n1281 ) : ( n1305 ) ;
assign n1307 =  ( n951 ) ? ( n1280 ) : ( n1306 ) ;
assign n1308 =  ( n950 ) ? ( n1279 ) : ( n1307 ) ;
assign n1309 =  ( n949 ) ? ( n1278 ) : ( n1308 ) ;
assign n1310 =  ( n947 ) ? ( n1277 ) : ( n1309 ) ;
assign n1311 =  ( n946 ) ? ( n1276 ) : ( n1310 ) ;
assign n1312 =  ( n943 ) ? ( n1275 ) : ( n1311 ) ;
assign n1313 =  ( n942 ) ? ( n1274 ) : ( n1312 ) ;
assign n1314 =  ( n939 ) ? ( n1273 ) : ( n1313 ) ;
assign n1315 =  ( n936 ) ? ( n1272 ) : ( n1314 ) ;
assign n1316 =  ( n934 ) ? ( n1271 ) : ( n1315 ) ;
assign n1317 =  ( n932 ) ? ( n1270 ) : ( n1316 ) ;
assign n1318 =  ( n930 ) ? ( n1269 ) : ( n1317 ) ;
assign n1319 =  ( n928 ) ? ( n1268 ) : ( n1318 ) ;
assign n1320 =  ( n926 ) ? ( n1267 ) : ( n1319 ) ;
assign n1321 =  ( n924 ) ? ( n1266 ) : ( n1320 ) ;
assign n1322 =  ( n621 ) ? ( n1321 ) : ( x12 ) ;
assign n1323 =  ( n1021 ) == ( 5'd13 )  ;
assign n1324 =  ( n1323 ) ? ( n1025 ) : ( x13 ) ;
assign n1325 =  ( n1323 ) ? ( n1027 ) : ( x13 ) ;
assign n1326 =  ( n1323 ) ? ( n1029 ) : ( x13 ) ;
assign n1327 =  ( n1323 ) ? ( n1031 ) : ( x13 ) ;
assign n1328 =  ( n1323 ) ? ( n1033 ) : ( x13 ) ;
assign n1329 =  ( n1323 ) ? ( n1035 ) : ( x13 ) ;
assign n1330 =  ( n1323 ) ? ( n1037 ) : ( x13 ) ;
assign n1331 =  ( n1323 ) ? ( n1039 ) : ( x13 ) ;
assign n1332 =  ( n1323 ) ? ( n1041 ) : ( x13 ) ;
assign n1333 =  ( n1323 ) ? ( n1043 ) : ( x13 ) ;
assign n1334 =  ( n1323 ) ? ( n1046 ) : ( x13 ) ;
assign n1335 =  ( n1323 ) ? ( n1048 ) : ( x13 ) ;
assign n1336 =  ( n1323 ) ? ( n1050 ) : ( x13 ) ;
assign n1337 =  ( n1323 ) ? ( n1053 ) : ( x13 ) ;
assign n1338 =  ( n1323 ) ? ( n1167 ) : ( x13 ) ;
assign n1339 =  ( n807 ) & ( n1055 )  ;
assign n1340 =  ( n1323 ) ? ( n1339 ) : ( x13 ) ;
assign n1341 =  ( n1323 ) ? ( n1283 ) : ( x13 ) ;
assign n1342 =  $signed( n807 ) < $signed( n1055 )  ;
assign n1343 =  ( n1342 ) ? ( 32'd1 ) : ( 32'd0 ) ;
assign n1344 =  ( n1323 ) ? ( n1343 ) : ( x13 ) ;
assign n1345 =  ( n1323 ) ? ( n1066 ) : ( x13 ) ;
assign n1346 =  ( n1323 ) ? ( n899 ) : ( x13 ) ;
assign n1347 =  ( n1323 ) ? ( n1072 ) : ( x13 ) ;
assign n1348 =  ( n1323 ) ? ( n1071 ) : ( x13 ) ;
assign n1349 =  ( n1323 ) ? ( n1097 ) : ( x13 ) ;
assign n1350 =  ( n1323 ) ? ( n1105 ) : ( x13 ) ;
assign n1351 =  ( n1323 ) ? ( n1114 ) : ( x13 ) ;
assign n1352 =  ( n1323 ) ? ( n1120 ) : ( x13 ) ;
assign n1353 =  ( n1323 ) ? ( n1122 ) : ( x13 ) ;
assign n1354 =  ( n967 ) ? ( n1353 ) : ( x13 ) ;
assign n1355 =  ( n966 ) ? ( n1352 ) : ( n1354 ) ;
assign n1356 =  ( n965 ) ? ( n1351 ) : ( n1355 ) ;
assign n1357 =  ( n964 ) ? ( n1350 ) : ( n1356 ) ;
assign n1358 =  ( n963 ) ? ( n1349 ) : ( n1357 ) ;
assign n1359 =  ( n957 ) ? ( n1348 ) : ( n1358 ) ;
assign n1360 =  ( n956 ) ? ( n1347 ) : ( n1359 ) ;
assign n1361 =  ( n1068 ) ? ( n1346 ) : ( n1360 ) ;
assign n1362 =  ( n955 ) ? ( n1345 ) : ( n1361 ) ;
assign n1363 =  ( n954 ) ? ( n1344 ) : ( n1362 ) ;
assign n1364 =  ( n953 ) ? ( n1341 ) : ( n1363 ) ;
assign n1365 =  ( n952 ) ? ( n1340 ) : ( n1364 ) ;
assign n1366 =  ( n951 ) ? ( n1338 ) : ( n1365 ) ;
assign n1367 =  ( n950 ) ? ( n1337 ) : ( n1366 ) ;
assign n1368 =  ( n949 ) ? ( n1336 ) : ( n1367 ) ;
assign n1369 =  ( n947 ) ? ( n1335 ) : ( n1368 ) ;
assign n1370 =  ( n946 ) ? ( n1334 ) : ( n1369 ) ;
assign n1371 =  ( n943 ) ? ( n1333 ) : ( n1370 ) ;
assign n1372 =  ( n942 ) ? ( n1332 ) : ( n1371 ) ;
assign n1373 =  ( n939 ) ? ( n1331 ) : ( n1372 ) ;
assign n1374 =  ( n936 ) ? ( n1330 ) : ( n1373 ) ;
assign n1375 =  ( n934 ) ? ( n1329 ) : ( n1374 ) ;
assign n1376 =  ( n932 ) ? ( n1328 ) : ( n1375 ) ;
assign n1377 =  ( n930 ) ? ( n1327 ) : ( n1376 ) ;
assign n1378 =  ( n928 ) ? ( n1326 ) : ( n1377 ) ;
assign n1379 =  ( n926 ) ? ( n1325 ) : ( n1378 ) ;
assign n1380 =  ( n924 ) ? ( n1324 ) : ( n1379 ) ;
assign n1381 =  ( n621 ) ? ( n1380 ) : ( x13 ) ;
assign n1382 =  ( n1021 ) == ( 5'd14 )  ;
assign n1383 =  ( n1382 ) ? ( n1025 ) : ( x14 ) ;
assign n1384 =  ( n1382 ) ? ( n1027 ) : ( x14 ) ;
assign n1385 =  ( n1382 ) ? ( n1029 ) : ( x14 ) ;
assign n1386 =  ( n1382 ) ? ( n1031 ) : ( x14 ) ;
assign n1387 =  ( n1382 ) ? ( n1033 ) : ( x14 ) ;
assign n1388 =  ( n1382 ) ? ( n1035 ) : ( x14 ) ;
assign n1389 =  ( n1382 ) ? ( n1037 ) : ( x14 ) ;
assign n1390 =  ( n1382 ) ? ( n1039 ) : ( x14 ) ;
assign n1391 =  ( n1382 ) ? ( n1041 ) : ( x14 ) ;
assign n1392 =  ( n1382 ) ? ( n1043 ) : ( x14 ) ;
assign n1393 =  ( n1382 ) ? ( n1046 ) : ( x14 ) ;
assign n1394 =  ( n1382 ) ? ( n1048 ) : ( x14 ) ;
assign n1395 =  ( n1382 ) ? ( n1050 ) : ( x14 ) ;
assign n1396 =  ( n1382 ) ? ( n1053 ) : ( x14 ) ;
assign n1397 =  ( n1382 ) ? ( n1167 ) : ( x14 ) ;
assign n1398 =  ( n1382 ) ? ( n1058 ) : ( x14 ) ;
assign n1399 =  ( n1382 ) ? ( n1283 ) : ( x14 ) ;
assign n1400 =  ( n1382 ) ? ( n1064 ) : ( x14 ) ;
assign n1401 =  ( n1382 ) ? ( n1066 ) : ( x14 ) ;
assign n1402 =  ( n1382 ) ? ( n899 ) : ( x14 ) ;
assign n1403 =  ( n1382 ) ? ( n1072 ) : ( x14 ) ;
assign n1404 =  ( n1382 ) ? ( n1071 ) : ( x14 ) ;
assign n1405 =  ( n1382 ) ? ( n1097 ) : ( x14 ) ;
assign n1406 =  ( n1382 ) ? ( n1105 ) : ( x14 ) ;
assign n1407 =  ( n1382 ) ? ( n1114 ) : ( x14 ) ;
assign n1408 =  ( n1382 ) ? ( n1120 ) : ( x14 ) ;
assign n1409 =  ( n1382 ) ? ( n1122 ) : ( x14 ) ;
assign n1410 =  ( n967 ) ? ( n1409 ) : ( x14 ) ;
assign n1411 =  ( n966 ) ? ( n1408 ) : ( n1410 ) ;
assign n1412 =  ( n965 ) ? ( n1407 ) : ( n1411 ) ;
assign n1413 =  ( n964 ) ? ( n1406 ) : ( n1412 ) ;
assign n1414 =  ( n963 ) ? ( n1405 ) : ( n1413 ) ;
assign n1415 =  ( n957 ) ? ( n1404 ) : ( n1414 ) ;
assign n1416 =  ( n956 ) ? ( n1403 ) : ( n1415 ) ;
assign n1417 =  ( n1068 ) ? ( n1402 ) : ( n1416 ) ;
assign n1418 =  ( n955 ) ? ( n1401 ) : ( n1417 ) ;
assign n1419 =  ( n954 ) ? ( n1400 ) : ( n1418 ) ;
assign n1420 =  ( n953 ) ? ( n1399 ) : ( n1419 ) ;
assign n1421 =  ( n952 ) ? ( n1398 ) : ( n1420 ) ;
assign n1422 =  ( n951 ) ? ( n1397 ) : ( n1421 ) ;
assign n1423 =  ( n950 ) ? ( n1396 ) : ( n1422 ) ;
assign n1424 =  ( n949 ) ? ( n1395 ) : ( n1423 ) ;
assign n1425 =  ( n947 ) ? ( n1394 ) : ( n1424 ) ;
assign n1426 =  ( n946 ) ? ( n1393 ) : ( n1425 ) ;
assign n1427 =  ( n943 ) ? ( n1392 ) : ( n1426 ) ;
assign n1428 =  ( n942 ) ? ( n1391 ) : ( n1427 ) ;
assign n1429 =  ( n939 ) ? ( n1390 ) : ( n1428 ) ;
assign n1430 =  ( n936 ) ? ( n1389 ) : ( n1429 ) ;
assign n1431 =  ( n934 ) ? ( n1388 ) : ( n1430 ) ;
assign n1432 =  ( n932 ) ? ( n1387 ) : ( n1431 ) ;
assign n1433 =  ( n930 ) ? ( n1386 ) : ( n1432 ) ;
assign n1434 =  ( n928 ) ? ( n1385 ) : ( n1433 ) ;
assign n1435 =  ( n926 ) ? ( n1384 ) : ( n1434 ) ;
assign n1436 =  ( n924 ) ? ( n1383 ) : ( n1435 ) ;
assign n1437 =  ( n621 ) ? ( n1436 ) : ( x14 ) ;
assign n1438 =  ( n1021 ) == ( 5'd15 )  ;
assign n1439 =  ( n1438 ) ? ( n1025 ) : ( x15 ) ;
assign n1440 =  ( n1438 ) ? ( n1027 ) : ( x15 ) ;
assign n1441 =  ( n1438 ) ? ( n1029 ) : ( x15 ) ;
assign n1442 =  ( n1438 ) ? ( n1031 ) : ( x15 ) ;
assign n1443 =  ( n1438 ) ? ( n1033 ) : ( x15 ) ;
assign n1444 =  ( n1438 ) ? ( n1035 ) : ( x15 ) ;
assign n1445 =  ( n1438 ) ? ( n1037 ) : ( x15 ) ;
assign n1446 =  ( n1438 ) ? ( n1039 ) : ( x15 ) ;
assign n1447 =  ( n1438 ) ? ( n1041 ) : ( x15 ) ;
assign n1448 =  ( n1438 ) ? ( n1043 ) : ( x15 ) ;
assign n1449 =  ( n1438 ) ? ( n1046 ) : ( x15 ) ;
assign n1450 =  ( n1438 ) ? ( n1048 ) : ( x15 ) ;
assign n1451 =  ( n1438 ) ? ( n1050 ) : ( x15 ) ;
assign n1452 =  ( n807 ) ^ ( n1055 )  ;
assign n1453 =  ( n1438 ) ? ( n1452 ) : ( x15 ) ;
assign n1454 =  ( n1438 ) ? ( n1167 ) : ( x15 ) ;
assign n1455 =  ( n1438 ) ? ( n1058 ) : ( x15 ) ;
assign n1456 =  ( n1438 ) ? ( n1061 ) : ( x15 ) ;
assign n1457 =  ( n1438 ) ? ( n1064 ) : ( x15 ) ;
assign n1458 =  ( n1438 ) ? ( n1066 ) : ( x15 ) ;
assign n1459 =  ( n1438 ) ? ( n899 ) : ( x15 ) ;
assign n1460 =  ( n1438 ) ? ( n1072 ) : ( x15 ) ;
assign n1461 =  ( n1438 ) ? ( n1071 ) : ( x15 ) ;
assign n1462 =  ( n1438 ) ? ( n1097 ) : ( x15 ) ;
assign n1463 =  ( n1438 ) ? ( n1105 ) : ( x15 ) ;
assign n1464 =  ( n1438 ) ? ( n1114 ) : ( x15 ) ;
assign n1465 =  ( n1438 ) ? ( n1120 ) : ( x15 ) ;
assign n1466 =  ( n1438 ) ? ( n1122 ) : ( x15 ) ;
assign n1467 =  ( n967 ) ? ( n1466 ) : ( x15 ) ;
assign n1468 =  ( n966 ) ? ( n1465 ) : ( n1467 ) ;
assign n1469 =  ( n965 ) ? ( n1464 ) : ( n1468 ) ;
assign n1470 =  ( n964 ) ? ( n1463 ) : ( n1469 ) ;
assign n1471 =  ( n963 ) ? ( n1462 ) : ( n1470 ) ;
assign n1472 =  ( n957 ) ? ( n1461 ) : ( n1471 ) ;
assign n1473 =  ( n956 ) ? ( n1460 ) : ( n1472 ) ;
assign n1474 =  ( n1068 ) ? ( n1459 ) : ( n1473 ) ;
assign n1475 =  ( n955 ) ? ( n1458 ) : ( n1474 ) ;
assign n1476 =  ( n954 ) ? ( n1457 ) : ( n1475 ) ;
assign n1477 =  ( n953 ) ? ( n1456 ) : ( n1476 ) ;
assign n1478 =  ( n952 ) ? ( n1455 ) : ( n1477 ) ;
assign n1479 =  ( n951 ) ? ( n1454 ) : ( n1478 ) ;
assign n1480 =  ( n950 ) ? ( n1453 ) : ( n1479 ) ;
assign n1481 =  ( n949 ) ? ( n1451 ) : ( n1480 ) ;
assign n1482 =  ( n947 ) ? ( n1450 ) : ( n1481 ) ;
assign n1483 =  ( n946 ) ? ( n1449 ) : ( n1482 ) ;
assign n1484 =  ( n943 ) ? ( n1448 ) : ( n1483 ) ;
assign n1485 =  ( n942 ) ? ( n1447 ) : ( n1484 ) ;
assign n1486 =  ( n939 ) ? ( n1446 ) : ( n1485 ) ;
assign n1487 =  ( n936 ) ? ( n1445 ) : ( n1486 ) ;
assign n1488 =  ( n934 ) ? ( n1444 ) : ( n1487 ) ;
assign n1489 =  ( n932 ) ? ( n1443 ) : ( n1488 ) ;
assign n1490 =  ( n930 ) ? ( n1442 ) : ( n1489 ) ;
assign n1491 =  ( n928 ) ? ( n1441 ) : ( n1490 ) ;
assign n1492 =  ( n926 ) ? ( n1440 ) : ( n1491 ) ;
assign n1493 =  ( n924 ) ? ( n1439 ) : ( n1492 ) ;
assign n1494 =  ( n621 ) ? ( n1493 ) : ( x15 ) ;
assign n1495 =  ( n1021 ) == ( 5'd16 )  ;
assign n1496 =  ( n1495 ) ? ( n1025 ) : ( x16 ) ;
assign n1497 =  ( n1495 ) ? ( n1027 ) : ( x16 ) ;
assign n1498 =  ( n1495 ) ? ( n1029 ) : ( x16 ) ;
assign n1499 =  ( n1495 ) ? ( n1031 ) : ( x16 ) ;
assign n1500 =  ( n1495 ) ? ( n1033 ) : ( x16 ) ;
assign n1501 =  ( n1495 ) ? ( n1035 ) : ( x16 ) ;
assign n1502 =  ( n1495 ) ? ( n1037 ) : ( x16 ) ;
assign n1503 =  ( n1495 ) ? ( n1039 ) : ( x16 ) ;
assign n1504 =  ( n1495 ) ? ( n1041 ) : ( x16 ) ;
assign n1505 =  ( n1495 ) ? ( n1043 ) : ( x16 ) ;
assign n1506 =  ( n1495 ) ? ( n1046 ) : ( x16 ) ;
assign n1507 =  ( n1495 ) ? ( n1048 ) : ( x16 ) ;
assign n1508 =  ( n1495 ) ? ( n1050 ) : ( x16 ) ;
assign n1509 =  ( n1495 ) ? ( n1053 ) : ( x16 ) ;
assign n1510 =  ( n1495 ) ? ( n1167 ) : ( x16 ) ;
assign n1511 =  ( n1495 ) ? ( n1058 ) : ( x16 ) ;
assign n1512 =  ( n1495 ) ? ( n1283 ) : ( x16 ) ;
assign n1513 =  ( n1495 ) ? ( n1064 ) : ( x16 ) ;
assign n1514 =  ( n1495 ) ? ( n1066 ) : ( x16 ) ;
assign n1515 =  ( n1495 ) ? ( n899 ) : ( x16 ) ;
assign n1516 =  ( n1495 ) ? ( n1072 ) : ( x16 ) ;
assign n1517 =  ( n1495 ) ? ( n1071 ) : ( x16 ) ;
assign n1518 =  ( n1495 ) ? ( n1097 ) : ( x16 ) ;
assign n1519 =  ( n1495 ) ? ( n1105 ) : ( x16 ) ;
assign n1520 =  ( n1495 ) ? ( n1114 ) : ( x16 ) ;
assign n1521 =  ( n1495 ) ? ( n1120 ) : ( x16 ) ;
assign n1522 =  ( n1495 ) ? ( n1122 ) : ( x16 ) ;
assign n1523 =  ( n967 ) ? ( n1522 ) : ( x16 ) ;
assign n1524 =  ( n966 ) ? ( n1521 ) : ( n1523 ) ;
assign n1525 =  ( n965 ) ? ( n1520 ) : ( n1524 ) ;
assign n1526 =  ( n964 ) ? ( n1519 ) : ( n1525 ) ;
assign n1527 =  ( n963 ) ? ( n1518 ) : ( n1526 ) ;
assign n1528 =  ( n957 ) ? ( n1517 ) : ( n1527 ) ;
assign n1529 =  ( n956 ) ? ( n1516 ) : ( n1528 ) ;
assign n1530 =  ( n1068 ) ? ( n1515 ) : ( n1529 ) ;
assign n1531 =  ( n955 ) ? ( n1514 ) : ( n1530 ) ;
assign n1532 =  ( n954 ) ? ( n1513 ) : ( n1531 ) ;
assign n1533 =  ( n953 ) ? ( n1512 ) : ( n1532 ) ;
assign n1534 =  ( n952 ) ? ( n1511 ) : ( n1533 ) ;
assign n1535 =  ( n951 ) ? ( n1510 ) : ( n1534 ) ;
assign n1536 =  ( n950 ) ? ( n1509 ) : ( n1535 ) ;
assign n1537 =  ( n949 ) ? ( n1508 ) : ( n1536 ) ;
assign n1538 =  ( n947 ) ? ( n1507 ) : ( n1537 ) ;
assign n1539 =  ( n946 ) ? ( n1506 ) : ( n1538 ) ;
assign n1540 =  ( n943 ) ? ( n1505 ) : ( n1539 ) ;
assign n1541 =  ( n942 ) ? ( n1504 ) : ( n1540 ) ;
assign n1542 =  ( n939 ) ? ( n1503 ) : ( n1541 ) ;
assign n1543 =  ( n936 ) ? ( n1502 ) : ( n1542 ) ;
assign n1544 =  ( n934 ) ? ( n1501 ) : ( n1543 ) ;
assign n1545 =  ( n932 ) ? ( n1500 ) : ( n1544 ) ;
assign n1546 =  ( n930 ) ? ( n1499 ) : ( n1545 ) ;
assign n1547 =  ( n928 ) ? ( n1498 ) : ( n1546 ) ;
assign n1548 =  ( n926 ) ? ( n1497 ) : ( n1547 ) ;
assign n1549 =  ( n924 ) ? ( n1496 ) : ( n1548 ) ;
assign n1550 =  ( n621 ) ? ( n1549 ) : ( x16 ) ;
assign n1551 =  ( n1021 ) == ( 5'd17 )  ;
assign n1552 =  ( n1551 ) ? ( n1025 ) : ( x17 ) ;
assign n1553 =  ( n1551 ) ? ( n1027 ) : ( x17 ) ;
assign n1554 =  ( n1551 ) ? ( n1029 ) : ( x17 ) ;
assign n1555 =  ( n1551 ) ? ( n1031 ) : ( x17 ) ;
assign n1556 =  ( n1551 ) ? ( n1033 ) : ( x17 ) ;
assign n1557 =  ( n1551 ) ? ( n1035 ) : ( x17 ) ;
assign n1558 =  ( n1551 ) ? ( n1037 ) : ( x17 ) ;
assign n1559 =  ( n1551 ) ? ( n1039 ) : ( x17 ) ;
assign n1560 =  ( n1551 ) ? ( n1041 ) : ( x17 ) ;
assign n1561 =  ( n1551 ) ? ( n1043 ) : ( x17 ) ;
assign n1562 =  ( n1551 ) ? ( n1046 ) : ( x17 ) ;
assign n1563 =  ( n1551 ) ? ( n1048 ) : ( x17 ) ;
assign n1564 =  ( n1551 ) ? ( n1050 ) : ( x17 ) ;
assign n1565 =  ( n1551 ) ? ( n1053 ) : ( x17 ) ;
assign n1566 =  ( n1551 ) ? ( n1167 ) : ( x17 ) ;
assign n1567 =  ( n1551 ) ? ( n1058 ) : ( x17 ) ;
assign n1568 =  ( n1551 ) ? ( n1283 ) : ( x17 ) ;
assign n1569 =  ( n1551 ) ? ( n1064 ) : ( x17 ) ;
assign n1570 =  ( n1551 ) ? ( n1066 ) : ( x17 ) ;
assign n1571 =  ( n1551 ) ? ( n899 ) : ( x17 ) ;
assign n1572 =  ( n1551 ) ? ( n1072 ) : ( x17 ) ;
assign n1573 =  ( n1551 ) ? ( n1071 ) : ( x17 ) ;
assign n1574 =  ( n1551 ) ? ( n1097 ) : ( x17 ) ;
assign n1575 =  ( n1551 ) ? ( n1105 ) : ( x17 ) ;
assign n1576 =  ( n1551 ) ? ( n1114 ) : ( x17 ) ;
assign n1577 =  ( n1551 ) ? ( n1120 ) : ( x17 ) ;
assign n1578 =  ( n1551 ) ? ( n1122 ) : ( x17 ) ;
assign n1579 =  ( n967 ) ? ( n1578 ) : ( x17 ) ;
assign n1580 =  ( n966 ) ? ( n1577 ) : ( n1579 ) ;
assign n1581 =  ( n965 ) ? ( n1576 ) : ( n1580 ) ;
assign n1582 =  ( n964 ) ? ( n1575 ) : ( n1581 ) ;
assign n1583 =  ( n963 ) ? ( n1574 ) : ( n1582 ) ;
assign n1584 =  ( n957 ) ? ( n1573 ) : ( n1583 ) ;
assign n1585 =  ( n956 ) ? ( n1572 ) : ( n1584 ) ;
assign n1586 =  ( n1068 ) ? ( n1571 ) : ( n1585 ) ;
assign n1587 =  ( n955 ) ? ( n1570 ) : ( n1586 ) ;
assign n1588 =  ( n954 ) ? ( n1569 ) : ( n1587 ) ;
assign n1589 =  ( n953 ) ? ( n1568 ) : ( n1588 ) ;
assign n1590 =  ( n952 ) ? ( n1567 ) : ( n1589 ) ;
assign n1591 =  ( n951 ) ? ( n1566 ) : ( n1590 ) ;
assign n1592 =  ( n950 ) ? ( n1565 ) : ( n1591 ) ;
assign n1593 =  ( n949 ) ? ( n1564 ) : ( n1592 ) ;
assign n1594 =  ( n947 ) ? ( n1563 ) : ( n1593 ) ;
assign n1595 =  ( n946 ) ? ( n1562 ) : ( n1594 ) ;
assign n1596 =  ( n943 ) ? ( n1561 ) : ( n1595 ) ;
assign n1597 =  ( n942 ) ? ( n1560 ) : ( n1596 ) ;
assign n1598 =  ( n939 ) ? ( n1559 ) : ( n1597 ) ;
assign n1599 =  ( n936 ) ? ( n1558 ) : ( n1598 ) ;
assign n1600 =  ( n934 ) ? ( n1557 ) : ( n1599 ) ;
assign n1601 =  ( n932 ) ? ( n1556 ) : ( n1600 ) ;
assign n1602 =  ( n930 ) ? ( n1555 ) : ( n1601 ) ;
assign n1603 =  ( n928 ) ? ( n1554 ) : ( n1602 ) ;
assign n1604 =  ( n926 ) ? ( n1553 ) : ( n1603 ) ;
assign n1605 =  ( n924 ) ? ( n1552 ) : ( n1604 ) ;
assign n1606 =  ( n621 ) ? ( n1605 ) : ( x17 ) ;
assign n1607 =  ( n1021 ) == ( 5'd18 )  ;
assign n1608 =  ( n1607 ) ? ( n1025 ) : ( x18 ) ;
assign n1609 =  ( n1607 ) ? ( n1027 ) : ( x18 ) ;
assign n1610 =  ( n1607 ) ? ( n1029 ) : ( x18 ) ;
assign n1611 =  ( n1607 ) ? ( n1031 ) : ( x18 ) ;
assign n1612 =  ( n1607 ) ? ( n1033 ) : ( x18 ) ;
assign n1613 =  ( n1607 ) ? ( n1035 ) : ( x18 ) ;
assign n1614 =  ( n1607 ) ? ( n1037 ) : ( x18 ) ;
assign n1615 =  ( n1607 ) ? ( n1039 ) : ( x18 ) ;
assign n1616 =  ( n1607 ) ? ( n1041 ) : ( x18 ) ;
assign n1617 =  ( n1607 ) ? ( n1043 ) : ( x18 ) ;
assign n1618 =  ( n1607 ) ? ( n1046 ) : ( x18 ) ;
assign n1619 =  ( n1607 ) ? ( n1048 ) : ( x18 ) ;
assign n1620 =  ( n1607 ) ? ( n1050 ) : ( x18 ) ;
assign n1621 =  ( n1607 ) ? ( n1053 ) : ( x18 ) ;
assign n1622 =  ( n1607 ) ? ( n1167 ) : ( x18 ) ;
assign n1623 =  ( n1607 ) ? ( n1339 ) : ( x18 ) ;
assign n1624 =  ( n1607 ) ? ( n1283 ) : ( x18 ) ;
assign n1625 =  ( n1607 ) ? ( n1064 ) : ( x18 ) ;
assign n1626 =  ( n1607 ) ? ( n1066 ) : ( x18 ) ;
assign n1627 =  ( n1607 ) ? ( n899 ) : ( x18 ) ;
assign n1628 =  ( n1607 ) ? ( n1072 ) : ( x18 ) ;
assign n1629 =  ( n1607 ) ? ( n1071 ) : ( x18 ) ;
assign n1630 =  ( n1607 ) ? ( n1097 ) : ( x18 ) ;
assign n1631 =  ( n1607 ) ? ( n1105 ) : ( x18 ) ;
assign n1632 =  ( n1607 ) ? ( n1114 ) : ( x18 ) ;
assign n1633 =  ( n1607 ) ? ( n1120 ) : ( x18 ) ;
assign n1634 =  ( n1607 ) ? ( n1122 ) : ( x18 ) ;
assign n1635 =  ( n967 ) ? ( n1634 ) : ( x18 ) ;
assign n1636 =  ( n966 ) ? ( n1633 ) : ( n1635 ) ;
assign n1637 =  ( n965 ) ? ( n1632 ) : ( n1636 ) ;
assign n1638 =  ( n964 ) ? ( n1631 ) : ( n1637 ) ;
assign n1639 =  ( n963 ) ? ( n1630 ) : ( n1638 ) ;
assign n1640 =  ( n957 ) ? ( n1629 ) : ( n1639 ) ;
assign n1641 =  ( n956 ) ? ( n1628 ) : ( n1640 ) ;
assign n1642 =  ( n1068 ) ? ( n1627 ) : ( n1641 ) ;
assign n1643 =  ( n955 ) ? ( n1626 ) : ( n1642 ) ;
assign n1644 =  ( n954 ) ? ( n1625 ) : ( n1643 ) ;
assign n1645 =  ( n953 ) ? ( n1624 ) : ( n1644 ) ;
assign n1646 =  ( n952 ) ? ( n1623 ) : ( n1645 ) ;
assign n1647 =  ( n951 ) ? ( n1622 ) : ( n1646 ) ;
assign n1648 =  ( n950 ) ? ( n1621 ) : ( n1647 ) ;
assign n1649 =  ( n949 ) ? ( n1620 ) : ( n1648 ) ;
assign n1650 =  ( n947 ) ? ( n1619 ) : ( n1649 ) ;
assign n1651 =  ( n946 ) ? ( n1618 ) : ( n1650 ) ;
assign n1652 =  ( n943 ) ? ( n1617 ) : ( n1651 ) ;
assign n1653 =  ( n942 ) ? ( n1616 ) : ( n1652 ) ;
assign n1654 =  ( n939 ) ? ( n1615 ) : ( n1653 ) ;
assign n1655 =  ( n936 ) ? ( n1614 ) : ( n1654 ) ;
assign n1656 =  ( n934 ) ? ( n1613 ) : ( n1655 ) ;
assign n1657 =  ( n932 ) ? ( n1612 ) : ( n1656 ) ;
assign n1658 =  ( n930 ) ? ( n1611 ) : ( n1657 ) ;
assign n1659 =  ( n928 ) ? ( n1610 ) : ( n1658 ) ;
assign n1660 =  ( n926 ) ? ( n1609 ) : ( n1659 ) ;
assign n1661 =  ( n924 ) ? ( n1608 ) : ( n1660 ) ;
assign n1662 =  ( n621 ) ? ( n1661 ) : ( x18 ) ;
assign n1663 =  ( n1021 ) == ( 5'd19 )  ;
assign n1664 =  ( n1663 ) ? ( n1025 ) : ( x19 ) ;
assign n1665 =  ( n1663 ) ? ( n1027 ) : ( x19 ) ;
assign n1666 =  ( n1663 ) ? ( n1029 ) : ( x19 ) ;
assign n1667 =  ( n1663 ) ? ( n1031 ) : ( x19 ) ;
assign n1668 =  ( n1663 ) ? ( n1033 ) : ( x19 ) ;
assign n1669 =  ( n1663 ) ? ( n1035 ) : ( x19 ) ;
assign n1670 =  ( n1663 ) ? ( n1037 ) : ( x19 ) ;
assign n1671 =  ( n1663 ) ? ( n1039 ) : ( x19 ) ;
assign n1672 =  ( n1663 ) ? ( n1041 ) : ( x19 ) ;
assign n1673 =  ( n1663 ) ? ( n1043 ) : ( x19 ) ;
assign n1674 =  ( n1663 ) ? ( n1046 ) : ( x19 ) ;
assign n1675 =  ( n1663 ) ? ( n1048 ) : ( x19 ) ;
assign n1676 =  ( n1663 ) ? ( n1050 ) : ( x19 ) ;
assign n1677 =  ( n1663 ) ? ( n1053 ) : ( x19 ) ;
assign n1678 =  ( n1663 ) ? ( n1056 ) : ( x19 ) ;
assign n1679 =  ( n1663 ) ? ( n1058 ) : ( x19 ) ;
assign n1680 =  ( n1663 ) ? ( n1283 ) : ( x19 ) ;
assign n1681 =  ( n1663 ) ? ( n1064 ) : ( x19 ) ;
assign n1682 =  ( n1663 ) ? ( n1066 ) : ( x19 ) ;
assign n1683 =  ( n1663 ) ? ( n899 ) : ( x19 ) ;
assign n1684 =  ( n1663 ) ? ( n1072 ) : ( x19 ) ;
assign n1685 =  ( n1663 ) ? ( n1071 ) : ( x19 ) ;
assign n1686 =  ( n1663 ) ? ( n1097 ) : ( x19 ) ;
assign n1687 =  ( n1663 ) ? ( n1105 ) : ( x19 ) ;
assign n1688 =  ( n1663 ) ? ( n1114 ) : ( x19 ) ;
assign n1689 =  ( n1663 ) ? ( n1120 ) : ( x19 ) ;
assign n1690 =  ( n1663 ) ? ( n1122 ) : ( x19 ) ;
assign n1691 =  ( n967 ) ? ( n1690 ) : ( x19 ) ;
assign n1692 =  ( n966 ) ? ( n1689 ) : ( n1691 ) ;
assign n1693 =  ( n965 ) ? ( n1688 ) : ( n1692 ) ;
assign n1694 =  ( n964 ) ? ( n1687 ) : ( n1693 ) ;
assign n1695 =  ( n963 ) ? ( n1686 ) : ( n1694 ) ;
assign n1696 =  ( n957 ) ? ( n1685 ) : ( n1695 ) ;
assign n1697 =  ( n956 ) ? ( n1684 ) : ( n1696 ) ;
assign n1698 =  ( n1068 ) ? ( n1683 ) : ( n1697 ) ;
assign n1699 =  ( n955 ) ? ( n1682 ) : ( n1698 ) ;
assign n1700 =  ( n954 ) ? ( n1681 ) : ( n1699 ) ;
assign n1701 =  ( n953 ) ? ( n1680 ) : ( n1700 ) ;
assign n1702 =  ( n952 ) ? ( n1679 ) : ( n1701 ) ;
assign n1703 =  ( n951 ) ? ( n1678 ) : ( n1702 ) ;
assign n1704 =  ( n950 ) ? ( n1677 ) : ( n1703 ) ;
assign n1705 =  ( n949 ) ? ( n1676 ) : ( n1704 ) ;
assign n1706 =  ( n947 ) ? ( n1675 ) : ( n1705 ) ;
assign n1707 =  ( n946 ) ? ( n1674 ) : ( n1706 ) ;
assign n1708 =  ( n943 ) ? ( n1673 ) : ( n1707 ) ;
assign n1709 =  ( n942 ) ? ( n1672 ) : ( n1708 ) ;
assign n1710 =  ( n939 ) ? ( n1671 ) : ( n1709 ) ;
assign n1711 =  ( n936 ) ? ( n1670 ) : ( n1710 ) ;
assign n1712 =  ( n934 ) ? ( n1669 ) : ( n1711 ) ;
assign n1713 =  ( n932 ) ? ( n1668 ) : ( n1712 ) ;
assign n1714 =  ( n930 ) ? ( n1667 ) : ( n1713 ) ;
assign n1715 =  ( n928 ) ? ( n1666 ) : ( n1714 ) ;
assign n1716 =  ( n926 ) ? ( n1665 ) : ( n1715 ) ;
assign n1717 =  ( n924 ) ? ( n1664 ) : ( n1716 ) ;
assign n1718 =  ( n621 ) ? ( n1717 ) : ( x19 ) ;
assign n1719 =  ( n1021 ) == ( 5'd2 )  ;
assign n1720 =  ( n1719 ) ? ( n1025 ) : ( x2 ) ;
assign n1721 =  ( n1719 ) ? ( n1027 ) : ( x2 ) ;
assign n1722 =  ( n1719 ) ? ( n1029 ) : ( x2 ) ;
assign n1723 =  ( n1719 ) ? ( n1031 ) : ( x2 ) ;
assign n1724 =  ( n1719 ) ? ( n1033 ) : ( x2 ) ;
assign n1725 =  ( n1719 ) ? ( n1035 ) : ( x2 ) ;
assign n1726 =  ( n1719 ) ? ( n1037 ) : ( x2 ) ;
assign n1727 =  ( n1719 ) ? ( n1039 ) : ( x2 ) ;
assign n1728 =  ( n1719 ) ? ( n1041 ) : ( x2 ) ;
assign n1729 =  ( n1719 ) ? ( n1043 ) : ( x2 ) ;
assign n1730 =  ( n1719 ) ? ( n1046 ) : ( x2 ) ;
assign n1731 =  ( n1719 ) ? ( n1048 ) : ( x2 ) ;
assign n1732 =  ( n1719 ) ? ( n1050 ) : ( x2 ) ;
assign n1733 =  ( n1719 ) ? ( n1053 ) : ( x2 ) ;
assign n1734 =  ( n1719 ) ? ( n1167 ) : ( x2 ) ;
assign n1735 =  ( n1719 ) ? ( n1058 ) : ( x2 ) ;
assign n1736 =  ( n1719 ) ? ( n1283 ) : ( x2 ) ;
assign n1737 =  ( n1719 ) ? ( n1064 ) : ( x2 ) ;
assign n1738 =  ( n1719 ) ? ( n1066 ) : ( x2 ) ;
assign n1739 =  ( n1719 ) ? ( n899 ) : ( x2 ) ;
assign n1740 =  ( n1719 ) ? ( n1072 ) : ( x2 ) ;
assign n1741 =  ( n1719 ) ? ( n1071 ) : ( x2 ) ;
assign n1742 =  ( n1719 ) ? ( n1097 ) : ( x2 ) ;
assign n1743 =  ( n1719 ) ? ( n1105 ) : ( x2 ) ;
assign n1744 =  ( n1719 ) ? ( n1114 ) : ( x2 ) ;
assign n1745 =  ( n1719 ) ? ( n1120 ) : ( x2 ) ;
assign n1746 =  ( n1719 ) ? ( n1122 ) : ( x2 ) ;
assign n1747 =  ( n967 ) ? ( n1746 ) : ( x2 ) ;
assign n1748 =  ( n966 ) ? ( n1745 ) : ( n1747 ) ;
assign n1749 =  ( n965 ) ? ( n1744 ) : ( n1748 ) ;
assign n1750 =  ( n964 ) ? ( n1743 ) : ( n1749 ) ;
assign n1751 =  ( n963 ) ? ( n1742 ) : ( n1750 ) ;
assign n1752 =  ( n957 ) ? ( n1741 ) : ( n1751 ) ;
assign n1753 =  ( n956 ) ? ( n1740 ) : ( n1752 ) ;
assign n1754 =  ( n1068 ) ? ( n1739 ) : ( n1753 ) ;
assign n1755 =  ( n955 ) ? ( n1738 ) : ( n1754 ) ;
assign n1756 =  ( n954 ) ? ( n1737 ) : ( n1755 ) ;
assign n1757 =  ( n953 ) ? ( n1736 ) : ( n1756 ) ;
assign n1758 =  ( n952 ) ? ( n1735 ) : ( n1757 ) ;
assign n1759 =  ( n951 ) ? ( n1734 ) : ( n1758 ) ;
assign n1760 =  ( n950 ) ? ( n1733 ) : ( n1759 ) ;
assign n1761 =  ( n949 ) ? ( n1732 ) : ( n1760 ) ;
assign n1762 =  ( n947 ) ? ( n1731 ) : ( n1761 ) ;
assign n1763 =  ( n946 ) ? ( n1730 ) : ( n1762 ) ;
assign n1764 =  ( n943 ) ? ( n1729 ) : ( n1763 ) ;
assign n1765 =  ( n942 ) ? ( n1728 ) : ( n1764 ) ;
assign n1766 =  ( n939 ) ? ( n1727 ) : ( n1765 ) ;
assign n1767 =  ( n936 ) ? ( n1726 ) : ( n1766 ) ;
assign n1768 =  ( n934 ) ? ( n1725 ) : ( n1767 ) ;
assign n1769 =  ( n932 ) ? ( n1724 ) : ( n1768 ) ;
assign n1770 =  ( n930 ) ? ( n1723 ) : ( n1769 ) ;
assign n1771 =  ( n928 ) ? ( n1722 ) : ( n1770 ) ;
assign n1772 =  ( n926 ) ? ( n1721 ) : ( n1771 ) ;
assign n1773 =  ( n924 ) ? ( n1720 ) : ( n1772 ) ;
assign n1774 =  ( n621 ) ? ( n1773 ) : ( x2 ) ;
assign n1775 =  ( n1021 ) == ( 5'd20 )  ;
assign n1776 =  ( n1775 ) ? ( n1025 ) : ( x20 ) ;
assign n1777 =  ( n1775 ) ? ( n1027 ) : ( x20 ) ;
assign n1778 =  ( n1775 ) ? ( n1029 ) : ( x20 ) ;
assign n1779 =  ( n1775 ) ? ( n1031 ) : ( x20 ) ;
assign n1780 =  ( n1775 ) ? ( n1033 ) : ( x20 ) ;
assign n1781 =  ( n1775 ) ? ( n1035 ) : ( x20 ) ;
assign n1782 =  ( n1775 ) ? ( n1037 ) : ( x20 ) ;
assign n1783 =  ( n1775 ) ? ( n1039 ) : ( x20 ) ;
assign n1784 =  ( n1775 ) ? ( n1041 ) : ( x20 ) ;
assign n1785 =  ( n1775 ) ? ( n1043 ) : ( x20 ) ;
assign n1786 =  ( n1775 ) ? ( n1046 ) : ( x20 ) ;
assign n1787 =  ( n1775 ) ? ( n1048 ) : ( x20 ) ;
assign n1788 =  ( n1775 ) ? ( n1050 ) : ( x20 ) ;
assign n1789 =  ( n1775 ) ? ( n1053 ) : ( x20 ) ;
assign n1790 =  ( n1775 ) ? ( n1167 ) : ( x20 ) ;
assign n1791 =  ( n1775 ) ? ( n1058 ) : ( x20 ) ;
assign n1792 =  ( n1775 ) ? ( n1061 ) : ( x20 ) ;
assign n1793 =  ( n1775 ) ? ( n1064 ) : ( x20 ) ;
assign n1794 =  ( n1775 ) ? ( n1066 ) : ( x20 ) ;
assign n1795 =  ( n1775 ) ? ( n899 ) : ( x20 ) ;
assign n1796 =  ( n1775 ) ? ( n1072 ) : ( x20 ) ;
assign n1797 =  ( n1775 ) ? ( n1071 ) : ( x20 ) ;
assign n1798 =  ( n1775 ) ? ( n1097 ) : ( x20 ) ;
assign n1799 =  ( n1775 ) ? ( n1105 ) : ( x20 ) ;
assign n1800 =  ( n1775 ) ? ( n1114 ) : ( x20 ) ;
assign n1801 =  ( n1775 ) ? ( n1120 ) : ( x20 ) ;
assign n1802 =  ( n1775 ) ? ( n1122 ) : ( x20 ) ;
assign n1803 =  ( n967 ) ? ( n1802 ) : ( x20 ) ;
assign n1804 =  ( n966 ) ? ( n1801 ) : ( n1803 ) ;
assign n1805 =  ( n965 ) ? ( n1800 ) : ( n1804 ) ;
assign n1806 =  ( n964 ) ? ( n1799 ) : ( n1805 ) ;
assign n1807 =  ( n963 ) ? ( n1798 ) : ( n1806 ) ;
assign n1808 =  ( n957 ) ? ( n1797 ) : ( n1807 ) ;
assign n1809 =  ( n956 ) ? ( n1796 ) : ( n1808 ) ;
assign n1810 =  ( n1068 ) ? ( n1795 ) : ( n1809 ) ;
assign n1811 =  ( n955 ) ? ( n1794 ) : ( n1810 ) ;
assign n1812 =  ( n954 ) ? ( n1793 ) : ( n1811 ) ;
assign n1813 =  ( n953 ) ? ( n1792 ) : ( n1812 ) ;
assign n1814 =  ( n952 ) ? ( n1791 ) : ( n1813 ) ;
assign n1815 =  ( n951 ) ? ( n1790 ) : ( n1814 ) ;
assign n1816 =  ( n950 ) ? ( n1789 ) : ( n1815 ) ;
assign n1817 =  ( n949 ) ? ( n1788 ) : ( n1816 ) ;
assign n1818 =  ( n947 ) ? ( n1787 ) : ( n1817 ) ;
assign n1819 =  ( n946 ) ? ( n1786 ) : ( n1818 ) ;
assign n1820 =  ( n943 ) ? ( n1785 ) : ( n1819 ) ;
assign n1821 =  ( n942 ) ? ( n1784 ) : ( n1820 ) ;
assign n1822 =  ( n939 ) ? ( n1783 ) : ( n1821 ) ;
assign n1823 =  ( n936 ) ? ( n1782 ) : ( n1822 ) ;
assign n1824 =  ( n934 ) ? ( n1781 ) : ( n1823 ) ;
assign n1825 =  ( n932 ) ? ( n1780 ) : ( n1824 ) ;
assign n1826 =  ( n930 ) ? ( n1779 ) : ( n1825 ) ;
assign n1827 =  ( n928 ) ? ( n1778 ) : ( n1826 ) ;
assign n1828 =  ( n926 ) ? ( n1777 ) : ( n1827 ) ;
assign n1829 =  ( n924 ) ? ( n1776 ) : ( n1828 ) ;
assign n1830 =  ( n621 ) ? ( n1829 ) : ( x20 ) ;
assign n1831 =  ( n1021 ) == ( 5'd21 )  ;
assign n1832 =  ( n1831 ) ? ( n1025 ) : ( x21 ) ;
assign n1833 =  ( n1831 ) ? ( n1027 ) : ( x21 ) ;
assign n1834 =  ( n1831 ) ? ( n1029 ) : ( x21 ) ;
assign n1835 =  ( n1831 ) ? ( n1031 ) : ( x21 ) ;
assign n1836 =  ( n1831 ) ? ( n1033 ) : ( x21 ) ;
assign n1837 =  ( n1831 ) ? ( n1035 ) : ( x21 ) ;
assign n1838 =  ( n1831 ) ? ( n1037 ) : ( x21 ) ;
assign n1839 =  ( n1831 ) ? ( n1039 ) : ( x21 ) ;
assign n1840 =  ( n1831 ) ? ( n1041 ) : ( x21 ) ;
assign n1841 =  ( n1831 ) ? ( n1043 ) : ( x21 ) ;
assign n1842 =  ( n1831 ) ? ( n1046 ) : ( x21 ) ;
assign n1843 =  ( n1831 ) ? ( n1048 ) : ( x21 ) ;
assign n1844 =  ( n1831 ) ? ( n1050 ) : ( x21 ) ;
assign n1845 =  ( n1831 ) ? ( n1053 ) : ( x21 ) ;
assign n1846 =  ( n1831 ) ? ( n1167 ) : ( x21 ) ;
assign n1847 =  ( n1831 ) ? ( n1339 ) : ( x21 ) ;
assign n1848 =  ( n1831 ) ? ( n1283 ) : ( x21 ) ;
assign n1849 =  ( n1831 ) ? ( n1343 ) : ( x21 ) ;
assign n1850 =  ( n1831 ) ? ( n1066 ) : ( x21 ) ;
assign n1851 =  ( n1831 ) ? ( n899 ) : ( x21 ) ;
assign n1852 =  ( n1831 ) ? ( n1072 ) : ( x21 ) ;
assign n1853 =  ( n1831 ) ? ( n1071 ) : ( x21 ) ;
assign n1854 =  ( n1831 ) ? ( n1097 ) : ( x21 ) ;
assign n1855 =  ( n1831 ) ? ( n1105 ) : ( x21 ) ;
assign n1856 =  ( n1831 ) ? ( n1114 ) : ( x21 ) ;
assign n1857 =  ( n1831 ) ? ( n1120 ) : ( x21 ) ;
assign n1858 =  ( n1831 ) ? ( n1122 ) : ( x21 ) ;
assign n1859 =  ( n967 ) ? ( n1858 ) : ( x21 ) ;
assign n1860 =  ( n966 ) ? ( n1857 ) : ( n1859 ) ;
assign n1861 =  ( n965 ) ? ( n1856 ) : ( n1860 ) ;
assign n1862 =  ( n964 ) ? ( n1855 ) : ( n1861 ) ;
assign n1863 =  ( n963 ) ? ( n1854 ) : ( n1862 ) ;
assign n1864 =  ( n957 ) ? ( n1853 ) : ( n1863 ) ;
assign n1865 =  ( n956 ) ? ( n1852 ) : ( n1864 ) ;
assign n1866 =  ( n1068 ) ? ( n1851 ) : ( n1865 ) ;
assign n1867 =  ( n955 ) ? ( n1850 ) : ( n1866 ) ;
assign n1868 =  ( n954 ) ? ( n1849 ) : ( n1867 ) ;
assign n1869 =  ( n953 ) ? ( n1848 ) : ( n1868 ) ;
assign n1870 =  ( n952 ) ? ( n1847 ) : ( n1869 ) ;
assign n1871 =  ( n951 ) ? ( n1846 ) : ( n1870 ) ;
assign n1872 =  ( n950 ) ? ( n1845 ) : ( n1871 ) ;
assign n1873 =  ( n949 ) ? ( n1844 ) : ( n1872 ) ;
assign n1874 =  ( n947 ) ? ( n1843 ) : ( n1873 ) ;
assign n1875 =  ( n946 ) ? ( n1842 ) : ( n1874 ) ;
assign n1876 =  ( n943 ) ? ( n1841 ) : ( n1875 ) ;
assign n1877 =  ( n942 ) ? ( n1840 ) : ( n1876 ) ;
assign n1878 =  ( n939 ) ? ( n1839 ) : ( n1877 ) ;
assign n1879 =  ( n936 ) ? ( n1838 ) : ( n1878 ) ;
assign n1880 =  ( n934 ) ? ( n1837 ) : ( n1879 ) ;
assign n1881 =  ( n932 ) ? ( n1836 ) : ( n1880 ) ;
assign n1882 =  ( n930 ) ? ( n1835 ) : ( n1881 ) ;
assign n1883 =  ( n928 ) ? ( n1834 ) : ( n1882 ) ;
assign n1884 =  ( n926 ) ? ( n1833 ) : ( n1883 ) ;
assign n1885 =  ( n924 ) ? ( n1832 ) : ( n1884 ) ;
assign n1886 =  ( n621 ) ? ( n1885 ) : ( x21 ) ;
assign n1887 =  ( n1021 ) == ( 5'd22 )  ;
assign n1888 =  ( n1887 ) ? ( n1025 ) : ( x22 ) ;
assign n1889 =  ( n1887 ) ? ( n1027 ) : ( x22 ) ;
assign n1890 =  ( n1887 ) ? ( n1029 ) : ( x22 ) ;
assign n1891 =  ( n1887 ) ? ( n1031 ) : ( x22 ) ;
assign n1892 =  ( n1887 ) ? ( n1033 ) : ( x22 ) ;
assign n1893 =  ( n1887 ) ? ( n1035 ) : ( x22 ) ;
assign n1894 =  ( n1887 ) ? ( n1037 ) : ( x22 ) ;
assign n1895 =  ( n1887 ) ? ( n1039 ) : ( x22 ) ;
assign n1896 =  ( n1887 ) ? ( n1041 ) : ( x22 ) ;
assign n1897 =  ( n1887 ) ? ( n1043 ) : ( x22 ) ;
assign n1898 =  ( n1887 ) ? ( n1046 ) : ( x22 ) ;
assign n1899 =  ( n1887 ) ? ( n1048 ) : ( x22 ) ;
assign n1900 =  ( n1887 ) ? ( n1050 ) : ( x22 ) ;
assign n1901 =  ( n1887 ) ? ( n1452 ) : ( x22 ) ;
assign n1902 =  ( n1887 ) ? ( n1167 ) : ( x22 ) ;
assign n1903 =  ( n1887 ) ? ( n1058 ) : ( x22 ) ;
assign n1904 =  ( n1887 ) ? ( n1061 ) : ( x22 ) ;
assign n1905 =  ( n1887 ) ? ( n1343 ) : ( x22 ) ;
assign n1906 =  ( n1887 ) ? ( n1066 ) : ( x22 ) ;
assign n1907 =  ( n1887 ) ? ( n899 ) : ( x22 ) ;
assign n1908 =  ( n1887 ) ? ( n1072 ) : ( x22 ) ;
assign n1909 =  ( n1887 ) ? ( n1071 ) : ( x22 ) ;
assign n1910 =  ( n1887 ) ? ( n1097 ) : ( x22 ) ;
assign n1911 =  ( n1887 ) ? ( n1105 ) : ( x22 ) ;
assign n1912 =  ( n1887 ) ? ( n1114 ) : ( x22 ) ;
assign n1913 =  ( n1887 ) ? ( n1120 ) : ( x22 ) ;
assign n1914 =  ( n1887 ) ? ( n1122 ) : ( x22 ) ;
assign n1915 =  ( n967 ) ? ( n1914 ) : ( x22 ) ;
assign n1916 =  ( n966 ) ? ( n1913 ) : ( n1915 ) ;
assign n1917 =  ( n965 ) ? ( n1912 ) : ( n1916 ) ;
assign n1918 =  ( n964 ) ? ( n1911 ) : ( n1917 ) ;
assign n1919 =  ( n963 ) ? ( n1910 ) : ( n1918 ) ;
assign n1920 =  ( n957 ) ? ( n1909 ) : ( n1919 ) ;
assign n1921 =  ( n956 ) ? ( n1908 ) : ( n1920 ) ;
assign n1922 =  ( n1068 ) ? ( n1907 ) : ( n1921 ) ;
assign n1923 =  ( n955 ) ? ( n1906 ) : ( n1922 ) ;
assign n1924 =  ( n954 ) ? ( n1905 ) : ( n1923 ) ;
assign n1925 =  ( n953 ) ? ( n1904 ) : ( n1924 ) ;
assign n1926 =  ( n952 ) ? ( n1903 ) : ( n1925 ) ;
assign n1927 =  ( n951 ) ? ( n1902 ) : ( n1926 ) ;
assign n1928 =  ( n950 ) ? ( n1901 ) : ( n1927 ) ;
assign n1929 =  ( n949 ) ? ( n1900 ) : ( n1928 ) ;
assign n1930 =  ( n947 ) ? ( n1899 ) : ( n1929 ) ;
assign n1931 =  ( n946 ) ? ( n1898 ) : ( n1930 ) ;
assign n1932 =  ( n943 ) ? ( n1897 ) : ( n1931 ) ;
assign n1933 =  ( n942 ) ? ( n1896 ) : ( n1932 ) ;
assign n1934 =  ( n939 ) ? ( n1895 ) : ( n1933 ) ;
assign n1935 =  ( n936 ) ? ( n1894 ) : ( n1934 ) ;
assign n1936 =  ( n934 ) ? ( n1893 ) : ( n1935 ) ;
assign n1937 =  ( n932 ) ? ( n1892 ) : ( n1936 ) ;
assign n1938 =  ( n930 ) ? ( n1891 ) : ( n1937 ) ;
assign n1939 =  ( n928 ) ? ( n1890 ) : ( n1938 ) ;
assign n1940 =  ( n926 ) ? ( n1889 ) : ( n1939 ) ;
assign n1941 =  ( n924 ) ? ( n1888 ) : ( n1940 ) ;
assign n1942 =  ( n621 ) ? ( n1941 ) : ( x22 ) ;
assign n1943 =  ( n1021 ) == ( 5'd23 )  ;
assign n1944 =  ( n1943 ) ? ( n1025 ) : ( x23 ) ;
assign n1945 =  ( n1943 ) ? ( n1027 ) : ( x23 ) ;
assign n1946 =  ( n1943 ) ? ( n1029 ) : ( x23 ) ;
assign n1947 =  ( n1943 ) ? ( n1031 ) : ( x23 ) ;
assign n1948 =  ( n1943 ) ? ( n1033 ) : ( x23 ) ;
assign n1949 =  ( n1943 ) ? ( n1035 ) : ( x23 ) ;
assign n1950 =  ( n1943 ) ? ( n1037 ) : ( x23 ) ;
assign n1951 =  ( n1943 ) ? ( n1039 ) : ( x23 ) ;
assign n1952 =  ( n1943 ) ? ( n1041 ) : ( x23 ) ;
assign n1953 =  ( n1943 ) ? ( n1043 ) : ( x23 ) ;
assign n1954 =  ( n1943 ) ? ( n1046 ) : ( x23 ) ;
assign n1955 =  ( n1943 ) ? ( n1048 ) : ( x23 ) ;
assign n1956 =  ( n1943 ) ? ( n1050 ) : ( x23 ) ;
assign n1957 =  ( n1943 ) ? ( n1452 ) : ( x23 ) ;
assign n1958 =  ( n1943 ) ? ( n1167 ) : ( x23 ) ;
assign n1959 =  ( n1943 ) ? ( n1058 ) : ( x23 ) ;
assign n1960 =  ( n1943 ) ? ( n1283 ) : ( x23 ) ;
assign n1961 =  ( n1943 ) ? ( n1343 ) : ( x23 ) ;
assign n1962 =  ( n1943 ) ? ( n1066 ) : ( x23 ) ;
assign n1963 =  ( n1943 ) ? ( n899 ) : ( x23 ) ;
assign n1964 =  ( n1943 ) ? ( n1072 ) : ( x23 ) ;
assign n1965 =  ( n1943 ) ? ( n1071 ) : ( x23 ) ;
assign n1966 =  ( n1943 ) ? ( n1097 ) : ( x23 ) ;
assign n1967 =  ( n1943 ) ? ( n1105 ) : ( x23 ) ;
assign n1968 =  ( n1943 ) ? ( n1114 ) : ( x23 ) ;
assign n1969 =  ( n1943 ) ? ( n1120 ) : ( x23 ) ;
assign n1970 =  ( n1943 ) ? ( n1122 ) : ( x23 ) ;
assign n1971 =  ( n967 ) ? ( n1970 ) : ( x23 ) ;
assign n1972 =  ( n966 ) ? ( n1969 ) : ( n1971 ) ;
assign n1973 =  ( n965 ) ? ( n1968 ) : ( n1972 ) ;
assign n1974 =  ( n964 ) ? ( n1967 ) : ( n1973 ) ;
assign n1975 =  ( n963 ) ? ( n1966 ) : ( n1974 ) ;
assign n1976 =  ( n957 ) ? ( n1965 ) : ( n1975 ) ;
assign n1977 =  ( n956 ) ? ( n1964 ) : ( n1976 ) ;
assign n1978 =  ( n1068 ) ? ( n1963 ) : ( n1977 ) ;
assign n1979 =  ( n955 ) ? ( n1962 ) : ( n1978 ) ;
assign n1980 =  ( n954 ) ? ( n1961 ) : ( n1979 ) ;
assign n1981 =  ( n953 ) ? ( n1960 ) : ( n1980 ) ;
assign n1982 =  ( n952 ) ? ( n1959 ) : ( n1981 ) ;
assign n1983 =  ( n951 ) ? ( n1958 ) : ( n1982 ) ;
assign n1984 =  ( n950 ) ? ( n1957 ) : ( n1983 ) ;
assign n1985 =  ( n949 ) ? ( n1956 ) : ( n1984 ) ;
assign n1986 =  ( n947 ) ? ( n1955 ) : ( n1985 ) ;
assign n1987 =  ( n946 ) ? ( n1954 ) : ( n1986 ) ;
assign n1988 =  ( n943 ) ? ( n1953 ) : ( n1987 ) ;
assign n1989 =  ( n942 ) ? ( n1952 ) : ( n1988 ) ;
assign n1990 =  ( n939 ) ? ( n1951 ) : ( n1989 ) ;
assign n1991 =  ( n936 ) ? ( n1950 ) : ( n1990 ) ;
assign n1992 =  ( n934 ) ? ( n1949 ) : ( n1991 ) ;
assign n1993 =  ( n932 ) ? ( n1948 ) : ( n1992 ) ;
assign n1994 =  ( n930 ) ? ( n1947 ) : ( n1993 ) ;
assign n1995 =  ( n928 ) ? ( n1946 ) : ( n1994 ) ;
assign n1996 =  ( n926 ) ? ( n1945 ) : ( n1995 ) ;
assign n1997 =  ( n924 ) ? ( n1944 ) : ( n1996 ) ;
assign n1998 =  ( n621 ) ? ( n1997 ) : ( x23 ) ;
assign n1999 =  ( n1021 ) == ( 5'd24 )  ;
assign n2000 =  ( n1999 ) ? ( n1025 ) : ( x24 ) ;
assign n2001 =  ( n1999 ) ? ( n1027 ) : ( x24 ) ;
assign n2002 =  ( n1999 ) ? ( n1029 ) : ( x24 ) ;
assign n2003 =  ( n1999 ) ? ( n1031 ) : ( x24 ) ;
assign n2004 =  ( n1999 ) ? ( n1033 ) : ( x24 ) ;
assign n2005 =  ( n1999 ) ? ( n1035 ) : ( x24 ) ;
assign n2006 =  ( n1999 ) ? ( n1037 ) : ( x24 ) ;
assign n2007 =  ( n1999 ) ? ( n1039 ) : ( x24 ) ;
assign n2008 =  ( n1999 ) ? ( n1041 ) : ( x24 ) ;
assign n2009 =  ( n1999 ) ? ( n1043 ) : ( x24 ) ;
assign n2010 =  ( n1999 ) ? ( n1046 ) : ( x24 ) ;
assign n2011 =  ( n1999 ) ? ( n1048 ) : ( x24 ) ;
assign n2012 =  ( n1999 ) ? ( n1050 ) : ( x24 ) ;
assign n2013 =  ( n1999 ) ? ( n1053 ) : ( x24 ) ;
assign n2014 =  ( n1999 ) ? ( n1167 ) : ( x24 ) ;
assign n2015 =  ( n1999 ) ? ( n1058 ) : ( x24 ) ;
assign n2016 =  ( n1999 ) ? ( n1283 ) : ( x24 ) ;
assign n2017 =  ( n1999 ) ? ( n1064 ) : ( x24 ) ;
assign n2018 =  ( n1999 ) ? ( n1066 ) : ( x24 ) ;
assign n2019 =  ( n1999 ) ? ( n899 ) : ( x24 ) ;
assign n2020 =  ( n1999 ) ? ( n1072 ) : ( x24 ) ;
assign n2021 =  ( n1999 ) ? ( n1071 ) : ( x24 ) ;
assign n2022 =  ( n1999 ) ? ( n1097 ) : ( x24 ) ;
assign n2023 =  ( n1999 ) ? ( n1105 ) : ( x24 ) ;
assign n2024 =  ( n1999 ) ? ( n1114 ) : ( x24 ) ;
assign n2025 =  ( n1999 ) ? ( n1120 ) : ( x24 ) ;
assign n2026 =  ( n1999 ) ? ( n1122 ) : ( x24 ) ;
assign n2027 =  ( n967 ) ? ( n2026 ) : ( x24 ) ;
assign n2028 =  ( n966 ) ? ( n2025 ) : ( n2027 ) ;
assign n2029 =  ( n965 ) ? ( n2024 ) : ( n2028 ) ;
assign n2030 =  ( n964 ) ? ( n2023 ) : ( n2029 ) ;
assign n2031 =  ( n963 ) ? ( n2022 ) : ( n2030 ) ;
assign n2032 =  ( n957 ) ? ( n2021 ) : ( n2031 ) ;
assign n2033 =  ( n956 ) ? ( n2020 ) : ( n2032 ) ;
assign n2034 =  ( n1068 ) ? ( n2019 ) : ( n2033 ) ;
assign n2035 =  ( n955 ) ? ( n2018 ) : ( n2034 ) ;
assign n2036 =  ( n954 ) ? ( n2017 ) : ( n2035 ) ;
assign n2037 =  ( n953 ) ? ( n2016 ) : ( n2036 ) ;
assign n2038 =  ( n952 ) ? ( n2015 ) : ( n2037 ) ;
assign n2039 =  ( n951 ) ? ( n2014 ) : ( n2038 ) ;
assign n2040 =  ( n950 ) ? ( n2013 ) : ( n2039 ) ;
assign n2041 =  ( n949 ) ? ( n2012 ) : ( n2040 ) ;
assign n2042 =  ( n947 ) ? ( n2011 ) : ( n2041 ) ;
assign n2043 =  ( n946 ) ? ( n2010 ) : ( n2042 ) ;
assign n2044 =  ( n943 ) ? ( n2009 ) : ( n2043 ) ;
assign n2045 =  ( n942 ) ? ( n2008 ) : ( n2044 ) ;
assign n2046 =  ( n939 ) ? ( n2007 ) : ( n2045 ) ;
assign n2047 =  ( n936 ) ? ( n2006 ) : ( n2046 ) ;
assign n2048 =  ( n934 ) ? ( n2005 ) : ( n2047 ) ;
assign n2049 =  ( n932 ) ? ( n2004 ) : ( n2048 ) ;
assign n2050 =  ( n930 ) ? ( n2003 ) : ( n2049 ) ;
assign n2051 =  ( n928 ) ? ( n2002 ) : ( n2050 ) ;
assign n2052 =  ( n926 ) ? ( n2001 ) : ( n2051 ) ;
assign n2053 =  ( n924 ) ? ( n2000 ) : ( n2052 ) ;
assign n2054 =  ( n621 ) ? ( n2053 ) : ( x24 ) ;
assign n2055 =  ( n1021 ) == ( 5'd25 )  ;
assign n2056 =  ( n2055 ) ? ( n1025 ) : ( x25 ) ;
assign n2057 =  ( n2055 ) ? ( n1027 ) : ( x25 ) ;
assign n2058 =  ( n2055 ) ? ( n1029 ) : ( x25 ) ;
assign n2059 =  ( n2055 ) ? ( n1031 ) : ( x25 ) ;
assign n2060 =  ( n2055 ) ? ( n1033 ) : ( x25 ) ;
assign n2061 =  ( n2055 ) ? ( n1035 ) : ( x25 ) ;
assign n2062 =  ( n2055 ) ? ( n1037 ) : ( x25 ) ;
assign n2063 =  ( n2055 ) ? ( n1039 ) : ( x25 ) ;
assign n2064 =  ( n2055 ) ? ( n1041 ) : ( x25 ) ;
assign n2065 =  ( n2055 ) ? ( n1043 ) : ( x25 ) ;
assign n2066 =  ( n2055 ) ? ( n1046 ) : ( x25 ) ;
assign n2067 =  ( n2055 ) ? ( n1048 ) : ( x25 ) ;
assign n2068 =  ( n2055 ) ? ( n1050 ) : ( x25 ) ;
assign n2069 =  ( n2055 ) ? ( n1053 ) : ( x25 ) ;
assign n2070 =  ( n2055 ) ? ( n1167 ) : ( x25 ) ;
assign n2071 =  ( n2055 ) ? ( n1058 ) : ( x25 ) ;
assign n2072 =  ( n2055 ) ? ( n1061 ) : ( x25 ) ;
assign n2073 =  ( n2055 ) ? ( n1064 ) : ( x25 ) ;
assign n2074 =  ( n2055 ) ? ( n1066 ) : ( x25 ) ;
assign n2075 =  ( n2055 ) ? ( n899 ) : ( x25 ) ;
assign n2076 =  ( n2055 ) ? ( n1072 ) : ( x25 ) ;
assign n2077 =  ( n2055 ) ? ( n1071 ) : ( x25 ) ;
assign n2078 =  ( n2055 ) ? ( n1097 ) : ( x25 ) ;
assign n2079 =  ( n2055 ) ? ( n1105 ) : ( x25 ) ;
assign n2080 =  ( n2055 ) ? ( n1114 ) : ( x25 ) ;
assign n2081 =  ( n2055 ) ? ( n1120 ) : ( x25 ) ;
assign n2082 =  ( n2055 ) ? ( n1122 ) : ( x25 ) ;
assign n2083 =  ( n967 ) ? ( n2082 ) : ( x25 ) ;
assign n2084 =  ( n966 ) ? ( n2081 ) : ( n2083 ) ;
assign n2085 =  ( n965 ) ? ( n2080 ) : ( n2084 ) ;
assign n2086 =  ( n964 ) ? ( n2079 ) : ( n2085 ) ;
assign n2087 =  ( n963 ) ? ( n2078 ) : ( n2086 ) ;
assign n2088 =  ( n957 ) ? ( n2077 ) : ( n2087 ) ;
assign n2089 =  ( n956 ) ? ( n2076 ) : ( n2088 ) ;
assign n2090 =  ( n1068 ) ? ( n2075 ) : ( n2089 ) ;
assign n2091 =  ( n955 ) ? ( n2074 ) : ( n2090 ) ;
assign n2092 =  ( n954 ) ? ( n2073 ) : ( n2091 ) ;
assign n2093 =  ( n953 ) ? ( n2072 ) : ( n2092 ) ;
assign n2094 =  ( n952 ) ? ( n2071 ) : ( n2093 ) ;
assign n2095 =  ( n951 ) ? ( n2070 ) : ( n2094 ) ;
assign n2096 =  ( n950 ) ? ( n2069 ) : ( n2095 ) ;
assign n2097 =  ( n949 ) ? ( n2068 ) : ( n2096 ) ;
assign n2098 =  ( n947 ) ? ( n2067 ) : ( n2097 ) ;
assign n2099 =  ( n946 ) ? ( n2066 ) : ( n2098 ) ;
assign n2100 =  ( n943 ) ? ( n2065 ) : ( n2099 ) ;
assign n2101 =  ( n942 ) ? ( n2064 ) : ( n2100 ) ;
assign n2102 =  ( n939 ) ? ( n2063 ) : ( n2101 ) ;
assign n2103 =  ( n936 ) ? ( n2062 ) : ( n2102 ) ;
assign n2104 =  ( n934 ) ? ( n2061 ) : ( n2103 ) ;
assign n2105 =  ( n932 ) ? ( n2060 ) : ( n2104 ) ;
assign n2106 =  ( n930 ) ? ( n2059 ) : ( n2105 ) ;
assign n2107 =  ( n928 ) ? ( n2058 ) : ( n2106 ) ;
assign n2108 =  ( n926 ) ? ( n2057 ) : ( n2107 ) ;
assign n2109 =  ( n924 ) ? ( n2056 ) : ( n2108 ) ;
assign n2110 =  ( n621 ) ? ( n2109 ) : ( x25 ) ;
assign n2111 =  ( n1021 ) == ( 5'd26 )  ;
assign n2112 =  ( n2111 ) ? ( n1025 ) : ( x26 ) ;
assign n2113 =  ( n2111 ) ? ( n1027 ) : ( x26 ) ;
assign n2114 =  ( n2111 ) ? ( n1029 ) : ( x26 ) ;
assign n2115 =  ( n2111 ) ? ( n1031 ) : ( x26 ) ;
assign n2116 =  ( n2111 ) ? ( n1033 ) : ( x26 ) ;
assign n2117 =  ( n2111 ) ? ( n1035 ) : ( x26 ) ;
assign n2118 =  ( n2111 ) ? ( n1037 ) : ( x26 ) ;
assign n2119 =  ( n2111 ) ? ( n1039 ) : ( x26 ) ;
assign n2120 =  ( n2111 ) ? ( n1041 ) : ( x26 ) ;
assign n2121 =  ( n2111 ) ? ( n1043 ) : ( x26 ) ;
assign n2122 =  ( n2111 ) ? ( n1046 ) : ( x26 ) ;
assign n2123 =  ( n2111 ) ? ( n1048 ) : ( x26 ) ;
assign n2124 =  ( n2111 ) ? ( n1050 ) : ( x26 ) ;
assign n2125 =  ( n2111 ) ? ( n1053 ) : ( x26 ) ;
assign n2126 =  ( n2111 ) ? ( n1167 ) : ( x26 ) ;
assign n2127 =  ( n2111 ) ? ( n1058 ) : ( x26 ) ;
assign n2128 =  ( n2111 ) ? ( n1283 ) : ( x26 ) ;
assign n2129 =  ( n2111 ) ? ( n1064 ) : ( x26 ) ;
assign n2130 =  ( n2111 ) ? ( n1066 ) : ( x26 ) ;
assign n2131 =  ( n2111 ) ? ( n899 ) : ( x26 ) ;
assign n2132 =  ( n2111 ) ? ( n1072 ) : ( x26 ) ;
assign n2133 =  ( n2111 ) ? ( n1071 ) : ( x26 ) ;
assign n2134 =  ( n2111 ) ? ( n1097 ) : ( x26 ) ;
assign n2135 =  ( n2111 ) ? ( n1105 ) : ( x26 ) ;
assign n2136 =  ( n2111 ) ? ( n1114 ) : ( x26 ) ;
assign n2137 =  ( n2111 ) ? ( n1120 ) : ( x26 ) ;
assign n2138 =  ( n2111 ) ? ( n1122 ) : ( x26 ) ;
assign n2139 =  ( n967 ) ? ( n2138 ) : ( x26 ) ;
assign n2140 =  ( n966 ) ? ( n2137 ) : ( n2139 ) ;
assign n2141 =  ( n965 ) ? ( n2136 ) : ( n2140 ) ;
assign n2142 =  ( n964 ) ? ( n2135 ) : ( n2141 ) ;
assign n2143 =  ( n963 ) ? ( n2134 ) : ( n2142 ) ;
assign n2144 =  ( n957 ) ? ( n2133 ) : ( n2143 ) ;
assign n2145 =  ( n956 ) ? ( n2132 ) : ( n2144 ) ;
assign n2146 =  ( n1068 ) ? ( n2131 ) : ( n2145 ) ;
assign n2147 =  ( n955 ) ? ( n2130 ) : ( n2146 ) ;
assign n2148 =  ( n954 ) ? ( n2129 ) : ( n2147 ) ;
assign n2149 =  ( n953 ) ? ( n2128 ) : ( n2148 ) ;
assign n2150 =  ( n952 ) ? ( n2127 ) : ( n2149 ) ;
assign n2151 =  ( n951 ) ? ( n2126 ) : ( n2150 ) ;
assign n2152 =  ( n950 ) ? ( n2125 ) : ( n2151 ) ;
assign n2153 =  ( n949 ) ? ( n2124 ) : ( n2152 ) ;
assign n2154 =  ( n947 ) ? ( n2123 ) : ( n2153 ) ;
assign n2155 =  ( n946 ) ? ( n2122 ) : ( n2154 ) ;
assign n2156 =  ( n943 ) ? ( n2121 ) : ( n2155 ) ;
assign n2157 =  ( n942 ) ? ( n2120 ) : ( n2156 ) ;
assign n2158 =  ( n939 ) ? ( n2119 ) : ( n2157 ) ;
assign n2159 =  ( n936 ) ? ( n2118 ) : ( n2158 ) ;
assign n2160 =  ( n934 ) ? ( n2117 ) : ( n2159 ) ;
assign n2161 =  ( n932 ) ? ( n2116 ) : ( n2160 ) ;
assign n2162 =  ( n930 ) ? ( n2115 ) : ( n2161 ) ;
assign n2163 =  ( n928 ) ? ( n2114 ) : ( n2162 ) ;
assign n2164 =  ( n926 ) ? ( n2113 ) : ( n2163 ) ;
assign n2165 =  ( n924 ) ? ( n2112 ) : ( n2164 ) ;
assign n2166 =  ( n621 ) ? ( n2165 ) : ( x26 ) ;
assign n2167 =  ( n1021 ) == ( 5'd27 )  ;
assign n2168 =  ( n2167 ) ? ( n1025 ) : ( x27 ) ;
assign n2169 =  ( n2167 ) ? ( n1027 ) : ( x27 ) ;
assign n2170 =  ( n2167 ) ? ( n1029 ) : ( x27 ) ;
assign n2171 =  ( n2167 ) ? ( n1031 ) : ( x27 ) ;
assign n2172 =  ( n2167 ) ? ( n1033 ) : ( x27 ) ;
assign n2173 =  ( n2167 ) ? ( n1035 ) : ( x27 ) ;
assign n2174 =  ( n2167 ) ? ( n1037 ) : ( x27 ) ;
assign n2175 =  ( n2167 ) ? ( n1039 ) : ( x27 ) ;
assign n2176 =  ( n2167 ) ? ( n1041 ) : ( x27 ) ;
assign n2177 =  ( n2167 ) ? ( n1043 ) : ( x27 ) ;
assign n2178 =  ( n2167 ) ? ( n1046 ) : ( x27 ) ;
assign n2179 =  ( n2167 ) ? ( n1048 ) : ( x27 ) ;
assign n2180 =  ( n2167 ) ? ( n1050 ) : ( x27 ) ;
assign n2181 =  ( n2167 ) ? ( n1053 ) : ( x27 ) ;
assign n2182 =  ( n2167 ) ? ( n1167 ) : ( x27 ) ;
assign n2183 =  ( n2167 ) ? ( n1339 ) : ( x27 ) ;
assign n2184 =  ( n2167 ) ? ( n1061 ) : ( x27 ) ;
assign n2185 =  ( n2167 ) ? ( n1064 ) : ( x27 ) ;
assign n2186 =  ( n2167 ) ? ( n1066 ) : ( x27 ) ;
assign n2187 =  ( n2167 ) ? ( n899 ) : ( x27 ) ;
assign n2188 =  ( n2167 ) ? ( n1072 ) : ( x27 ) ;
assign n2189 =  ( n2167 ) ? ( n1071 ) : ( x27 ) ;
assign n2190 =  ( n2167 ) ? ( n1097 ) : ( x27 ) ;
assign n2191 =  ( n2167 ) ? ( n1105 ) : ( x27 ) ;
assign n2192 =  ( n2167 ) ? ( n1114 ) : ( x27 ) ;
assign n2193 =  ( n2167 ) ? ( n1120 ) : ( x27 ) ;
assign n2194 =  ( n2167 ) ? ( n1122 ) : ( x27 ) ;
assign n2195 =  ( n967 ) ? ( n2194 ) : ( x27 ) ;
assign n2196 =  ( n966 ) ? ( n2193 ) : ( n2195 ) ;
assign n2197 =  ( n965 ) ? ( n2192 ) : ( n2196 ) ;
assign n2198 =  ( n964 ) ? ( n2191 ) : ( n2197 ) ;
assign n2199 =  ( n963 ) ? ( n2190 ) : ( n2198 ) ;
assign n2200 =  ( n957 ) ? ( n2189 ) : ( n2199 ) ;
assign n2201 =  ( n956 ) ? ( n2188 ) : ( n2200 ) ;
assign n2202 =  ( n1068 ) ? ( n2187 ) : ( n2201 ) ;
assign n2203 =  ( n955 ) ? ( n2186 ) : ( n2202 ) ;
assign n2204 =  ( n954 ) ? ( n2185 ) : ( n2203 ) ;
assign n2205 =  ( n953 ) ? ( n2184 ) : ( n2204 ) ;
assign n2206 =  ( n952 ) ? ( n2183 ) : ( n2205 ) ;
assign n2207 =  ( n951 ) ? ( n2182 ) : ( n2206 ) ;
assign n2208 =  ( n950 ) ? ( n2181 ) : ( n2207 ) ;
assign n2209 =  ( n949 ) ? ( n2180 ) : ( n2208 ) ;
assign n2210 =  ( n947 ) ? ( n2179 ) : ( n2209 ) ;
assign n2211 =  ( n946 ) ? ( n2178 ) : ( n2210 ) ;
assign n2212 =  ( n943 ) ? ( n2177 ) : ( n2211 ) ;
assign n2213 =  ( n942 ) ? ( n2176 ) : ( n2212 ) ;
assign n2214 =  ( n939 ) ? ( n2175 ) : ( n2213 ) ;
assign n2215 =  ( n936 ) ? ( n2174 ) : ( n2214 ) ;
assign n2216 =  ( n934 ) ? ( n2173 ) : ( n2215 ) ;
assign n2217 =  ( n932 ) ? ( n2172 ) : ( n2216 ) ;
assign n2218 =  ( n930 ) ? ( n2171 ) : ( n2217 ) ;
assign n2219 =  ( n928 ) ? ( n2170 ) : ( n2218 ) ;
assign n2220 =  ( n926 ) ? ( n2169 ) : ( n2219 ) ;
assign n2221 =  ( n924 ) ? ( n2168 ) : ( n2220 ) ;
assign n2222 =  ( n621 ) ? ( n2221 ) : ( x27 ) ;
assign n2223 =  ( n1021 ) == ( 5'd28 )  ;
assign n2224 =  ( n2223 ) ? ( n1025 ) : ( x28 ) ;
assign n2225 =  ( n2223 ) ? ( n1027 ) : ( x28 ) ;
assign n2226 =  ( n2223 ) ? ( n1029 ) : ( x28 ) ;
assign n2227 =  ( n2223 ) ? ( n1031 ) : ( x28 ) ;
assign n2228 =  ( n2223 ) ? ( n1033 ) : ( x28 ) ;
assign n2229 =  ( n2223 ) ? ( n1035 ) : ( x28 ) ;
assign n2230 =  ( n2223 ) ? ( n1037 ) : ( x28 ) ;
assign n2231 =  ( n2223 ) ? ( n1039 ) : ( x28 ) ;
assign n2232 =  ( n2223 ) ? ( n1041 ) : ( x28 ) ;
assign n2233 =  ( n2223 ) ? ( n1043 ) : ( x28 ) ;
assign n2234 =  ( n2223 ) ? ( n1046 ) : ( x28 ) ;
assign n2235 =  ( n2223 ) ? ( n1048 ) : ( x28 ) ;
assign n2236 =  ( n2223 ) ? ( n1050 ) : ( x28 ) ;
assign n2237 =  ( n2223 ) ? ( n1053 ) : ( x28 ) ;
assign n2238 =  ( n2223 ) ? ( n1167 ) : ( x28 ) ;
assign n2239 =  ( n2223 ) ? ( n1058 ) : ( x28 ) ;
assign n2240 =  ( n2223 ) ? ( n1061 ) : ( x28 ) ;
assign n2241 =  ( n2223 ) ? ( n1064 ) : ( x28 ) ;
assign n2242 =  ( n2223 ) ? ( n1066 ) : ( x28 ) ;
assign n2243 =  ( n2223 ) ? ( n899 ) : ( x28 ) ;
assign n2244 =  ( n2223 ) ? ( n1072 ) : ( x28 ) ;
assign n2245 =  ( n2223 ) ? ( n1071 ) : ( x28 ) ;
assign n2246 =  ( n2223 ) ? ( n1097 ) : ( x28 ) ;
assign n2247 =  ( n2223 ) ? ( n1105 ) : ( x28 ) ;
assign n2248 =  ( n2223 ) ? ( n1114 ) : ( x28 ) ;
assign n2249 =  ( n2223 ) ? ( n1120 ) : ( x28 ) ;
assign n2250 =  ( n2223 ) ? ( n1122 ) : ( x28 ) ;
assign n2251 =  ( n967 ) ? ( n2250 ) : ( x28 ) ;
assign n2252 =  ( n966 ) ? ( n2249 ) : ( n2251 ) ;
assign n2253 =  ( n965 ) ? ( n2248 ) : ( n2252 ) ;
assign n2254 =  ( n964 ) ? ( n2247 ) : ( n2253 ) ;
assign n2255 =  ( n963 ) ? ( n2246 ) : ( n2254 ) ;
assign n2256 =  ( n957 ) ? ( n2245 ) : ( n2255 ) ;
assign n2257 =  ( n956 ) ? ( n2244 ) : ( n2256 ) ;
assign n2258 =  ( n1068 ) ? ( n2243 ) : ( n2257 ) ;
assign n2259 =  ( n955 ) ? ( n2242 ) : ( n2258 ) ;
assign n2260 =  ( n954 ) ? ( n2241 ) : ( n2259 ) ;
assign n2261 =  ( n953 ) ? ( n2240 ) : ( n2260 ) ;
assign n2262 =  ( n952 ) ? ( n2239 ) : ( n2261 ) ;
assign n2263 =  ( n951 ) ? ( n2238 ) : ( n2262 ) ;
assign n2264 =  ( n950 ) ? ( n2237 ) : ( n2263 ) ;
assign n2265 =  ( n949 ) ? ( n2236 ) : ( n2264 ) ;
assign n2266 =  ( n947 ) ? ( n2235 ) : ( n2265 ) ;
assign n2267 =  ( n946 ) ? ( n2234 ) : ( n2266 ) ;
assign n2268 =  ( n943 ) ? ( n2233 ) : ( n2267 ) ;
assign n2269 =  ( n942 ) ? ( n2232 ) : ( n2268 ) ;
assign n2270 =  ( n939 ) ? ( n2231 ) : ( n2269 ) ;
assign n2271 =  ( n936 ) ? ( n2230 ) : ( n2270 ) ;
assign n2272 =  ( n934 ) ? ( n2229 ) : ( n2271 ) ;
assign n2273 =  ( n932 ) ? ( n2228 ) : ( n2272 ) ;
assign n2274 =  ( n930 ) ? ( n2227 ) : ( n2273 ) ;
assign n2275 =  ( n928 ) ? ( n2226 ) : ( n2274 ) ;
assign n2276 =  ( n926 ) ? ( n2225 ) : ( n2275 ) ;
assign n2277 =  ( n924 ) ? ( n2224 ) : ( n2276 ) ;
assign n2278 =  ( n621 ) ? ( n2277 ) : ( x28 ) ;
assign n2279 =  ( n1021 ) == ( 5'd29 )  ;
assign n2280 =  ( n2279 ) ? ( n1025 ) : ( x29 ) ;
assign n2281 =  ( n2279 ) ? ( n1027 ) : ( x29 ) ;
assign n2282 =  ( n2279 ) ? ( n1029 ) : ( x29 ) ;
assign n2283 =  ( n2279 ) ? ( n1031 ) : ( x29 ) ;
assign n2284 =  ( n2279 ) ? ( n1033 ) : ( x29 ) ;
assign n2285 =  ( n2279 ) ? ( n1035 ) : ( x29 ) ;
assign n2286 =  ( n2279 ) ? ( n1037 ) : ( x29 ) ;
assign n2287 =  ( n2279 ) ? ( n1039 ) : ( x29 ) ;
assign n2288 =  ( n2279 ) ? ( n1041 ) : ( x29 ) ;
assign n2289 =  ( n2279 ) ? ( n1043 ) : ( x29 ) ;
assign n2290 =  ( n2279 ) ? ( n1046 ) : ( x29 ) ;
assign n2291 =  ( n2279 ) ? ( n1048 ) : ( x29 ) ;
assign n2292 =  ( n2279 ) ? ( n1050 ) : ( x29 ) ;
assign n2293 =  ( n2279 ) ? ( n1053 ) : ( x29 ) ;
assign n2294 =  ( n2279 ) ? ( n1167 ) : ( x29 ) ;
assign n2295 =  ( n2279 ) ? ( n1339 ) : ( x29 ) ;
assign n2296 =  ( n2279 ) ? ( n1283 ) : ( x29 ) ;
assign n2297 =  ( n2279 ) ? ( n1343 ) : ( x29 ) ;
assign n2298 =  ( n2279 ) ? ( n1066 ) : ( x29 ) ;
assign n2299 =  ( n2279 ) ? ( n899 ) : ( x29 ) ;
assign n2300 =  ( n2279 ) ? ( n1072 ) : ( x29 ) ;
assign n2301 =  ( n2279 ) ? ( n1071 ) : ( x29 ) ;
assign n2302 =  ( n2279 ) ? ( n1097 ) : ( x29 ) ;
assign n2303 =  ( n2279 ) ? ( n1105 ) : ( x29 ) ;
assign n2304 =  ( n2279 ) ? ( n1114 ) : ( x29 ) ;
assign n2305 =  ( n2279 ) ? ( n1120 ) : ( x29 ) ;
assign n2306 =  ( n2279 ) ? ( n1122 ) : ( x29 ) ;
assign n2307 =  ( n967 ) ? ( n2306 ) : ( x29 ) ;
assign n2308 =  ( n966 ) ? ( n2305 ) : ( n2307 ) ;
assign n2309 =  ( n965 ) ? ( n2304 ) : ( n2308 ) ;
assign n2310 =  ( n964 ) ? ( n2303 ) : ( n2309 ) ;
assign n2311 =  ( n963 ) ? ( n2302 ) : ( n2310 ) ;
assign n2312 =  ( n957 ) ? ( n2301 ) : ( n2311 ) ;
assign n2313 =  ( n956 ) ? ( n2300 ) : ( n2312 ) ;
assign n2314 =  ( n1068 ) ? ( n2299 ) : ( n2313 ) ;
assign n2315 =  ( n955 ) ? ( n2298 ) : ( n2314 ) ;
assign n2316 =  ( n954 ) ? ( n2297 ) : ( n2315 ) ;
assign n2317 =  ( n953 ) ? ( n2296 ) : ( n2316 ) ;
assign n2318 =  ( n952 ) ? ( n2295 ) : ( n2317 ) ;
assign n2319 =  ( n951 ) ? ( n2294 ) : ( n2318 ) ;
assign n2320 =  ( n950 ) ? ( n2293 ) : ( n2319 ) ;
assign n2321 =  ( n949 ) ? ( n2292 ) : ( n2320 ) ;
assign n2322 =  ( n947 ) ? ( n2291 ) : ( n2321 ) ;
assign n2323 =  ( n946 ) ? ( n2290 ) : ( n2322 ) ;
assign n2324 =  ( n943 ) ? ( n2289 ) : ( n2323 ) ;
assign n2325 =  ( n942 ) ? ( n2288 ) : ( n2324 ) ;
assign n2326 =  ( n939 ) ? ( n2287 ) : ( n2325 ) ;
assign n2327 =  ( n936 ) ? ( n2286 ) : ( n2326 ) ;
assign n2328 =  ( n934 ) ? ( n2285 ) : ( n2327 ) ;
assign n2329 =  ( n932 ) ? ( n2284 ) : ( n2328 ) ;
assign n2330 =  ( n930 ) ? ( n2283 ) : ( n2329 ) ;
assign n2331 =  ( n928 ) ? ( n2282 ) : ( n2330 ) ;
assign n2332 =  ( n926 ) ? ( n2281 ) : ( n2331 ) ;
assign n2333 =  ( n924 ) ? ( n2280 ) : ( n2332 ) ;
assign n2334 =  ( n621 ) ? ( n2333 ) : ( x29 ) ;
assign n2335 =  ( n1021 ) == ( 5'd3 )  ;
assign n2336 =  ( n2335 ) ? ( n1025 ) : ( x3 ) ;
assign n2337 =  ( n2335 ) ? ( n1027 ) : ( x3 ) ;
assign n2338 =  ( n2335 ) ? ( n1029 ) : ( x3 ) ;
assign n2339 =  ( n2335 ) ? ( n1031 ) : ( x3 ) ;
assign n2340 =  ( n2335 ) ? ( n1033 ) : ( x3 ) ;
assign n2341 =  ( n2335 ) ? ( n1035 ) : ( x3 ) ;
assign n2342 =  ( n2335 ) ? ( n1037 ) : ( x3 ) ;
assign n2343 =  ( n2335 ) ? ( n1039 ) : ( x3 ) ;
assign n2344 =  ( n2335 ) ? ( n1041 ) : ( x3 ) ;
assign n2345 =  ( n2335 ) ? ( n1043 ) : ( x3 ) ;
assign n2346 =  ( n2335 ) ? ( n1046 ) : ( x3 ) ;
assign n2347 =  ( n2335 ) ? ( n1048 ) : ( x3 ) ;
assign n2348 =  ( n2335 ) ? ( n1050 ) : ( x3 ) ;
assign n2349 =  ( n2335 ) ? ( n1053 ) : ( x3 ) ;
assign n2350 =  ( n2335 ) ? ( n1167 ) : ( x3 ) ;
assign n2351 =  ( n2335 ) ? ( n1339 ) : ( x3 ) ;
assign n2352 =  ( n2335 ) ? ( n1061 ) : ( x3 ) ;
assign n2353 =  ( n2335 ) ? ( n1064 ) : ( x3 ) ;
assign n2354 =  ( n2335 ) ? ( n1066 ) : ( x3 ) ;
assign n2355 =  ( n2335 ) ? ( n899 ) : ( x3 ) ;
assign n2356 =  ( n2335 ) ? ( n1072 ) : ( x3 ) ;
assign n2357 =  ( n2335 ) ? ( n1071 ) : ( x3 ) ;
assign n2358 =  ( n2335 ) ? ( n1097 ) : ( x3 ) ;
assign n2359 =  ( n2335 ) ? ( n1105 ) : ( x3 ) ;
assign n2360 =  ( n2335 ) ? ( n1114 ) : ( x3 ) ;
assign n2361 =  ( n2335 ) ? ( n1120 ) : ( x3 ) ;
assign n2362 =  ( n2335 ) ? ( n1122 ) : ( x3 ) ;
assign n2363 =  ( n967 ) ? ( n2362 ) : ( x3 ) ;
assign n2364 =  ( n966 ) ? ( n2361 ) : ( n2363 ) ;
assign n2365 =  ( n965 ) ? ( n2360 ) : ( n2364 ) ;
assign n2366 =  ( n964 ) ? ( n2359 ) : ( n2365 ) ;
assign n2367 =  ( n963 ) ? ( n2358 ) : ( n2366 ) ;
assign n2368 =  ( n957 ) ? ( n2357 ) : ( n2367 ) ;
assign n2369 =  ( n956 ) ? ( n2356 ) : ( n2368 ) ;
assign n2370 =  ( n1068 ) ? ( n2355 ) : ( n2369 ) ;
assign n2371 =  ( n955 ) ? ( n2354 ) : ( n2370 ) ;
assign n2372 =  ( n954 ) ? ( n2353 ) : ( n2371 ) ;
assign n2373 =  ( n953 ) ? ( n2352 ) : ( n2372 ) ;
assign n2374 =  ( n952 ) ? ( n2351 ) : ( n2373 ) ;
assign n2375 =  ( n951 ) ? ( n2350 ) : ( n2374 ) ;
assign n2376 =  ( n950 ) ? ( n2349 ) : ( n2375 ) ;
assign n2377 =  ( n949 ) ? ( n2348 ) : ( n2376 ) ;
assign n2378 =  ( n947 ) ? ( n2347 ) : ( n2377 ) ;
assign n2379 =  ( n946 ) ? ( n2346 ) : ( n2378 ) ;
assign n2380 =  ( n943 ) ? ( n2345 ) : ( n2379 ) ;
assign n2381 =  ( n942 ) ? ( n2344 ) : ( n2380 ) ;
assign n2382 =  ( n939 ) ? ( n2343 ) : ( n2381 ) ;
assign n2383 =  ( n936 ) ? ( n2342 ) : ( n2382 ) ;
assign n2384 =  ( n934 ) ? ( n2341 ) : ( n2383 ) ;
assign n2385 =  ( n932 ) ? ( n2340 ) : ( n2384 ) ;
assign n2386 =  ( n930 ) ? ( n2339 ) : ( n2385 ) ;
assign n2387 =  ( n928 ) ? ( n2338 ) : ( n2386 ) ;
assign n2388 =  ( n926 ) ? ( n2337 ) : ( n2387 ) ;
assign n2389 =  ( n924 ) ? ( n2336 ) : ( n2388 ) ;
assign n2390 =  ( n621 ) ? ( n2389 ) : ( x3 ) ;
assign n2391 =  ( n1021 ) == ( 5'd30 )  ;
assign n2392 =  ( n2391 ) ? ( n1025 ) : ( x30 ) ;
assign n2393 =  ( n2391 ) ? ( n1027 ) : ( x30 ) ;
assign n2394 =  ( n2391 ) ? ( n1029 ) : ( x30 ) ;
assign n2395 =  ( n2391 ) ? ( n1031 ) : ( x30 ) ;
assign n2396 =  ( n2391 ) ? ( n1033 ) : ( x30 ) ;
assign n2397 =  ( n2391 ) ? ( n1035 ) : ( x30 ) ;
assign n2398 =  ( n2391 ) ? ( n1037 ) : ( x30 ) ;
assign n2399 =  ( n2391 ) ? ( n1039 ) : ( x30 ) ;
assign n2400 =  ( n2391 ) ? ( n1041 ) : ( x30 ) ;
assign n2401 =  ( n2391 ) ? ( n1043 ) : ( x30 ) ;
assign n2402 =  ( n2391 ) ? ( n1046 ) : ( x30 ) ;
assign n2403 =  ( n2391 ) ? ( n1048 ) : ( x30 ) ;
assign n2404 =  ( n2391 ) ? ( n1050 ) : ( x30 ) ;
assign n2405 =  ( n2391 ) ? ( n1053 ) : ( x30 ) ;
assign n2406 =  ( n2391 ) ? ( n1167 ) : ( x30 ) ;
assign n2407 =  ( n2391 ) ? ( n1058 ) : ( x30 ) ;
assign n2408 =  ( n2391 ) ? ( n1283 ) : ( x30 ) ;
assign n2409 =  ( n2391 ) ? ( n1064 ) : ( x30 ) ;
assign n2410 =  ( n2391 ) ? ( n1066 ) : ( x30 ) ;
assign n2411 =  ( n2391 ) ? ( n899 ) : ( x30 ) ;
assign n2412 =  ( n2391 ) ? ( n1072 ) : ( x30 ) ;
assign n2413 =  ( n2391 ) ? ( n1071 ) : ( x30 ) ;
assign n2414 =  ( n2391 ) ? ( n1097 ) : ( x30 ) ;
assign n2415 =  ( n2391 ) ? ( n1105 ) : ( x30 ) ;
assign n2416 =  ( n2391 ) ? ( n1114 ) : ( x30 ) ;
assign n2417 =  ( n2391 ) ? ( n1120 ) : ( x30 ) ;
assign n2418 =  ( n2391 ) ? ( n1122 ) : ( x30 ) ;
assign n2419 =  ( n967 ) ? ( n2418 ) : ( x30 ) ;
assign n2420 =  ( n966 ) ? ( n2417 ) : ( n2419 ) ;
assign n2421 =  ( n965 ) ? ( n2416 ) : ( n2420 ) ;
assign n2422 =  ( n964 ) ? ( n2415 ) : ( n2421 ) ;
assign n2423 =  ( n963 ) ? ( n2414 ) : ( n2422 ) ;
assign n2424 =  ( n957 ) ? ( n2413 ) : ( n2423 ) ;
assign n2425 =  ( n956 ) ? ( n2412 ) : ( n2424 ) ;
assign n2426 =  ( n1068 ) ? ( n2411 ) : ( n2425 ) ;
assign n2427 =  ( n955 ) ? ( n2410 ) : ( n2426 ) ;
assign n2428 =  ( n954 ) ? ( n2409 ) : ( n2427 ) ;
assign n2429 =  ( n953 ) ? ( n2408 ) : ( n2428 ) ;
assign n2430 =  ( n952 ) ? ( n2407 ) : ( n2429 ) ;
assign n2431 =  ( n951 ) ? ( n2406 ) : ( n2430 ) ;
assign n2432 =  ( n950 ) ? ( n2405 ) : ( n2431 ) ;
assign n2433 =  ( n949 ) ? ( n2404 ) : ( n2432 ) ;
assign n2434 =  ( n947 ) ? ( n2403 ) : ( n2433 ) ;
assign n2435 =  ( n946 ) ? ( n2402 ) : ( n2434 ) ;
assign n2436 =  ( n943 ) ? ( n2401 ) : ( n2435 ) ;
assign n2437 =  ( n942 ) ? ( n2400 ) : ( n2436 ) ;
assign n2438 =  ( n939 ) ? ( n2399 ) : ( n2437 ) ;
assign n2439 =  ( n936 ) ? ( n2398 ) : ( n2438 ) ;
assign n2440 =  ( n934 ) ? ( n2397 ) : ( n2439 ) ;
assign n2441 =  ( n932 ) ? ( n2396 ) : ( n2440 ) ;
assign n2442 =  ( n930 ) ? ( n2395 ) : ( n2441 ) ;
assign n2443 =  ( n928 ) ? ( n2394 ) : ( n2442 ) ;
assign n2444 =  ( n926 ) ? ( n2393 ) : ( n2443 ) ;
assign n2445 =  ( n924 ) ? ( n2392 ) : ( n2444 ) ;
assign n2446 =  ( n621 ) ? ( n2445 ) : ( x30 ) ;
assign n2447 =  ( n1021 ) == ( 5'd31 )  ;
assign n2448 =  ( n2447 ) ? ( n1025 ) : ( x31 ) ;
assign n2449 =  ( n2447 ) ? ( n1027 ) : ( x31 ) ;
assign n2450 =  ( n2447 ) ? ( n1029 ) : ( x31 ) ;
assign n2451 =  ( n2447 ) ? ( n1031 ) : ( x31 ) ;
assign n2452 =  ( n2447 ) ? ( n1033 ) : ( x31 ) ;
assign n2453 =  ( n2447 ) ? ( n1035 ) : ( x31 ) ;
assign n2454 =  ( n2447 ) ? ( n1037 ) : ( x31 ) ;
assign n2455 =  ( n2447 ) ? ( n1039 ) : ( x31 ) ;
assign n2456 =  ( n2447 ) ? ( n1041 ) : ( x31 ) ;
assign n2457 =  ( n2447 ) ? ( n1043 ) : ( x31 ) ;
assign n2458 =  ( n2447 ) ? ( n1046 ) : ( x31 ) ;
assign n2459 =  ( n2447 ) ? ( n1048 ) : ( x31 ) ;
assign n2460 =  ( n2447 ) ? ( n1050 ) : ( x31 ) ;
assign n2461 =  ( n2447 ) ? ( n1053 ) : ( x31 ) ;
assign n2462 =  ( n2447 ) ? ( n1167 ) : ( x31 ) ;
assign n2463 =  ( n2447 ) ? ( n1058 ) : ( x31 ) ;
assign n2464 =  ( n2447 ) ? ( n1283 ) : ( x31 ) ;
assign n2465 =  ( n2447 ) ? ( n1064 ) : ( x31 ) ;
assign n2466 =  ( n2447 ) ? ( n1066 ) : ( x31 ) ;
assign n2467 =  ( n2447 ) ? ( n899 ) : ( x31 ) ;
assign n2468 =  ( n2447 ) ? ( n1072 ) : ( x31 ) ;
assign n2469 =  ( n2447 ) ? ( n1071 ) : ( x31 ) ;
assign n2470 =  ( n2447 ) ? ( n1097 ) : ( x31 ) ;
assign n2471 =  ( n2447 ) ? ( n1105 ) : ( x31 ) ;
assign n2472 =  ( n2447 ) ? ( n1114 ) : ( x31 ) ;
assign n2473 =  ( n2447 ) ? ( n1120 ) : ( x31 ) ;
assign n2474 =  ( n2447 ) ? ( n1122 ) : ( x31 ) ;
assign n2475 =  ( n967 ) ? ( n2474 ) : ( x31 ) ;
assign n2476 =  ( n966 ) ? ( n2473 ) : ( n2475 ) ;
assign n2477 =  ( n965 ) ? ( n2472 ) : ( n2476 ) ;
assign n2478 =  ( n964 ) ? ( n2471 ) : ( n2477 ) ;
assign n2479 =  ( n963 ) ? ( n2470 ) : ( n2478 ) ;
assign n2480 =  ( n957 ) ? ( n2469 ) : ( n2479 ) ;
assign n2481 =  ( n956 ) ? ( n2468 ) : ( n2480 ) ;
assign n2482 =  ( n1068 ) ? ( n2467 ) : ( n2481 ) ;
assign n2483 =  ( n955 ) ? ( n2466 ) : ( n2482 ) ;
assign n2484 =  ( n954 ) ? ( n2465 ) : ( n2483 ) ;
assign n2485 =  ( n953 ) ? ( n2464 ) : ( n2484 ) ;
assign n2486 =  ( n952 ) ? ( n2463 ) : ( n2485 ) ;
assign n2487 =  ( n951 ) ? ( n2462 ) : ( n2486 ) ;
assign n2488 =  ( n950 ) ? ( n2461 ) : ( n2487 ) ;
assign n2489 =  ( n949 ) ? ( n2460 ) : ( n2488 ) ;
assign n2490 =  ( n947 ) ? ( n2459 ) : ( n2489 ) ;
assign n2491 =  ( n946 ) ? ( n2458 ) : ( n2490 ) ;
assign n2492 =  ( n943 ) ? ( n2457 ) : ( n2491 ) ;
assign n2493 =  ( n942 ) ? ( n2456 ) : ( n2492 ) ;
assign n2494 =  ( n939 ) ? ( n2455 ) : ( n2493 ) ;
assign n2495 =  ( n936 ) ? ( n2454 ) : ( n2494 ) ;
assign n2496 =  ( n934 ) ? ( n2453 ) : ( n2495 ) ;
assign n2497 =  ( n932 ) ? ( n2452 ) : ( n2496 ) ;
assign n2498 =  ( n930 ) ? ( n2451 ) : ( n2497 ) ;
assign n2499 =  ( n928 ) ? ( n2450 ) : ( n2498 ) ;
assign n2500 =  ( n926 ) ? ( n2449 ) : ( n2499 ) ;
assign n2501 =  ( n924 ) ? ( n2448 ) : ( n2500 ) ;
assign n2502 =  ( n621 ) ? ( n2501 ) : ( x31 ) ;
assign n2503 =  ( n1021 ) == ( 5'd4 )  ;
assign n2504 =  ( n2503 ) ? ( n1025 ) : ( x4 ) ;
assign n2505 =  ( n2503 ) ? ( n1027 ) : ( x4 ) ;
assign n2506 =  ( n2503 ) ? ( n1029 ) : ( x4 ) ;
assign n2507 =  ( n2503 ) ? ( n1031 ) : ( x4 ) ;
assign n2508 =  ( n2503 ) ? ( n1033 ) : ( x4 ) ;
assign n2509 =  ( n2503 ) ? ( n1035 ) : ( x4 ) ;
assign n2510 =  ( n2503 ) ? ( n1037 ) : ( x4 ) ;
assign n2511 =  ( n2503 ) ? ( n1039 ) : ( x4 ) ;
assign n2512 =  ( n2503 ) ? ( n1041 ) : ( x4 ) ;
assign n2513 =  ( n2503 ) ? ( n1043 ) : ( x4 ) ;
assign n2514 =  ( n2503 ) ? ( n1046 ) : ( x4 ) ;
assign n2515 =  ( n2503 ) ? ( n1048 ) : ( x4 ) ;
assign n2516 =  ( n2503 ) ? ( n1050 ) : ( x4 ) ;
assign n2517 =  ( n2503 ) ? ( n1053 ) : ( x4 ) ;
assign n2518 =  ( n2503 ) ? ( n1167 ) : ( x4 ) ;
assign n2519 =  ( n2503 ) ? ( n1058 ) : ( x4 ) ;
assign n2520 =  ( n2503 ) ? ( n1283 ) : ( x4 ) ;
assign n2521 =  ( n2503 ) ? ( n1064 ) : ( x4 ) ;
assign n2522 =  ( n2503 ) ? ( n1066 ) : ( x4 ) ;
assign n2523 =  ( n2503 ) ? ( n899 ) : ( x4 ) ;
assign n2524 =  ( n2503 ) ? ( n1072 ) : ( x4 ) ;
assign n2525 =  ( n2503 ) ? ( n1071 ) : ( x4 ) ;
assign n2526 =  ( n2503 ) ? ( n1097 ) : ( x4 ) ;
assign n2527 =  ( n2503 ) ? ( n1105 ) : ( x4 ) ;
assign n2528 =  ( n2503 ) ? ( n1114 ) : ( x4 ) ;
assign n2529 =  ( n2503 ) ? ( n1120 ) : ( x4 ) ;
assign n2530 =  ( n2503 ) ? ( n1122 ) : ( x4 ) ;
assign n2531 =  ( n967 ) ? ( n2530 ) : ( x4 ) ;
assign n2532 =  ( n966 ) ? ( n2529 ) : ( n2531 ) ;
assign n2533 =  ( n965 ) ? ( n2528 ) : ( n2532 ) ;
assign n2534 =  ( n964 ) ? ( n2527 ) : ( n2533 ) ;
assign n2535 =  ( n963 ) ? ( n2526 ) : ( n2534 ) ;
assign n2536 =  ( n957 ) ? ( n2525 ) : ( n2535 ) ;
assign n2537 =  ( n956 ) ? ( n2524 ) : ( n2536 ) ;
assign n2538 =  ( n1068 ) ? ( n2523 ) : ( n2537 ) ;
assign n2539 =  ( n955 ) ? ( n2522 ) : ( n2538 ) ;
assign n2540 =  ( n954 ) ? ( n2521 ) : ( n2539 ) ;
assign n2541 =  ( n953 ) ? ( n2520 ) : ( n2540 ) ;
assign n2542 =  ( n952 ) ? ( n2519 ) : ( n2541 ) ;
assign n2543 =  ( n951 ) ? ( n2518 ) : ( n2542 ) ;
assign n2544 =  ( n950 ) ? ( n2517 ) : ( n2543 ) ;
assign n2545 =  ( n949 ) ? ( n2516 ) : ( n2544 ) ;
assign n2546 =  ( n947 ) ? ( n2515 ) : ( n2545 ) ;
assign n2547 =  ( n946 ) ? ( n2514 ) : ( n2546 ) ;
assign n2548 =  ( n943 ) ? ( n2513 ) : ( n2547 ) ;
assign n2549 =  ( n942 ) ? ( n2512 ) : ( n2548 ) ;
assign n2550 =  ( n939 ) ? ( n2511 ) : ( n2549 ) ;
assign n2551 =  ( n936 ) ? ( n2510 ) : ( n2550 ) ;
assign n2552 =  ( n934 ) ? ( n2509 ) : ( n2551 ) ;
assign n2553 =  ( n932 ) ? ( n2508 ) : ( n2552 ) ;
assign n2554 =  ( n930 ) ? ( n2507 ) : ( n2553 ) ;
assign n2555 =  ( n928 ) ? ( n2506 ) : ( n2554 ) ;
assign n2556 =  ( n926 ) ? ( n2505 ) : ( n2555 ) ;
assign n2557 =  ( n924 ) ? ( n2504 ) : ( n2556 ) ;
assign n2558 =  ( n621 ) ? ( n2557 ) : ( x4 ) ;
assign n2559 =  ( n1021 ) == ( 5'd5 )  ;
assign n2560 =  ( n2559 ) ? ( n1025 ) : ( x5 ) ;
assign n2561 =  ( n2559 ) ? ( n1027 ) : ( x5 ) ;
assign n2562 =  ( n2559 ) ? ( n1029 ) : ( x5 ) ;
assign n2563 =  ( n2559 ) ? ( n1031 ) : ( x5 ) ;
assign n2564 =  ( n2559 ) ? ( n1033 ) : ( x5 ) ;
assign n2565 =  ( n2559 ) ? ( n1035 ) : ( x5 ) ;
assign n2566 =  ( n2559 ) ? ( n1037 ) : ( x5 ) ;
assign n2567 =  ( n2559 ) ? ( n1039 ) : ( x5 ) ;
assign n2568 =  ( n2559 ) ? ( n1041 ) : ( x5 ) ;
assign n2569 =  ( n2559 ) ? ( n1043 ) : ( x5 ) ;
assign n2570 =  ( n2559 ) ? ( n1046 ) : ( x5 ) ;
assign n2571 =  ( n2559 ) ? ( n1048 ) : ( x5 ) ;
assign n2572 =  ( n2559 ) ? ( n1050 ) : ( x5 ) ;
assign n2573 =  ( n2559 ) ? ( n1053 ) : ( x5 ) ;
assign n2574 =  ( n2559 ) ? ( n1167 ) : ( x5 ) ;
assign n2575 =  ( n2559 ) ? ( n1058 ) : ( x5 ) ;
assign n2576 =  ( n2559 ) ? ( n1061 ) : ( x5 ) ;
assign n2577 =  ( n2559 ) ? ( n1343 ) : ( x5 ) ;
assign n2578 =  ( n2559 ) ? ( n1066 ) : ( x5 ) ;
assign n2579 =  ( n2559 ) ? ( n899 ) : ( x5 ) ;
assign n2580 =  ( n2559 ) ? ( n1072 ) : ( x5 ) ;
assign n2581 =  ( n2559 ) ? ( n1071 ) : ( x5 ) ;
assign n2582 =  ( n2559 ) ? ( n1097 ) : ( x5 ) ;
assign n2583 =  ( n2559 ) ? ( n1105 ) : ( x5 ) ;
assign n2584 =  ( n2559 ) ? ( n1114 ) : ( x5 ) ;
assign n2585 =  ( n2559 ) ? ( n1120 ) : ( x5 ) ;
assign n2586 =  ( n2559 ) ? ( n1122 ) : ( x5 ) ;
assign n2587 =  ( n967 ) ? ( n2586 ) : ( x5 ) ;
assign n2588 =  ( n966 ) ? ( n2585 ) : ( n2587 ) ;
assign n2589 =  ( n965 ) ? ( n2584 ) : ( n2588 ) ;
assign n2590 =  ( n964 ) ? ( n2583 ) : ( n2589 ) ;
assign n2591 =  ( n963 ) ? ( n2582 ) : ( n2590 ) ;
assign n2592 =  ( n957 ) ? ( n2581 ) : ( n2591 ) ;
assign n2593 =  ( n956 ) ? ( n2580 ) : ( n2592 ) ;
assign n2594 =  ( n1068 ) ? ( n2579 ) : ( n2593 ) ;
assign n2595 =  ( n955 ) ? ( n2578 ) : ( n2594 ) ;
assign n2596 =  ( n954 ) ? ( n2577 ) : ( n2595 ) ;
assign n2597 =  ( n953 ) ? ( n2576 ) : ( n2596 ) ;
assign n2598 =  ( n952 ) ? ( n2575 ) : ( n2597 ) ;
assign n2599 =  ( n951 ) ? ( n2574 ) : ( n2598 ) ;
assign n2600 =  ( n950 ) ? ( n2573 ) : ( n2599 ) ;
assign n2601 =  ( n949 ) ? ( n2572 ) : ( n2600 ) ;
assign n2602 =  ( n947 ) ? ( n2571 ) : ( n2601 ) ;
assign n2603 =  ( n946 ) ? ( n2570 ) : ( n2602 ) ;
assign n2604 =  ( n943 ) ? ( n2569 ) : ( n2603 ) ;
assign n2605 =  ( n942 ) ? ( n2568 ) : ( n2604 ) ;
assign n2606 =  ( n939 ) ? ( n2567 ) : ( n2605 ) ;
assign n2607 =  ( n936 ) ? ( n2566 ) : ( n2606 ) ;
assign n2608 =  ( n934 ) ? ( n2565 ) : ( n2607 ) ;
assign n2609 =  ( n932 ) ? ( n2564 ) : ( n2608 ) ;
assign n2610 =  ( n930 ) ? ( n2563 ) : ( n2609 ) ;
assign n2611 =  ( n928 ) ? ( n2562 ) : ( n2610 ) ;
assign n2612 =  ( n926 ) ? ( n2561 ) : ( n2611 ) ;
assign n2613 =  ( n924 ) ? ( n2560 ) : ( n2612 ) ;
assign n2614 =  ( n621 ) ? ( n2613 ) : ( x5 ) ;
assign n2615 =  ( n1021 ) == ( 5'd6 )  ;
assign n2616 =  ( n2615 ) ? ( n1025 ) : ( x6 ) ;
assign n2617 =  ( n2615 ) ? ( n1027 ) : ( x6 ) ;
assign n2618 =  ( n2615 ) ? ( n1029 ) : ( x6 ) ;
assign n2619 =  ( n2615 ) ? ( n1031 ) : ( x6 ) ;
assign n2620 =  ( n2615 ) ? ( n1033 ) : ( x6 ) ;
assign n2621 =  ( n2615 ) ? ( n1035 ) : ( x6 ) ;
assign n2622 =  ( n2615 ) ? ( n1037 ) : ( x6 ) ;
assign n2623 =  ( n2615 ) ? ( n1039 ) : ( x6 ) ;
assign n2624 =  ( n2615 ) ? ( n1041 ) : ( x6 ) ;
assign n2625 =  ( n2615 ) ? ( n1043 ) : ( x6 ) ;
assign n2626 =  ( n2615 ) ? ( n1046 ) : ( x6 ) ;
assign n2627 =  ( n2615 ) ? ( n1048 ) : ( x6 ) ;
assign n2628 =  ( n2615 ) ? ( n1050 ) : ( x6 ) ;
assign n2629 =  ( n2615 ) ? ( n1053 ) : ( x6 ) ;
assign n2630 =  ( n2615 ) ? ( n1167 ) : ( x6 ) ;
assign n2631 =  ( n2615 ) ? ( n1058 ) : ( x6 ) ;
assign n2632 =  ( n2615 ) ? ( n1283 ) : ( x6 ) ;
assign n2633 =  ( n2615 ) ? ( n1064 ) : ( x6 ) ;
assign n2634 =  ( n807 ) + ( n1055 )  ;
assign n2635 =  ( n2615 ) ? ( n2634 ) : ( x6 ) ;
assign n2636 =  ( n2615 ) ? ( n899 ) : ( x6 ) ;
assign n2637 =  ( n2615 ) ? ( n1072 ) : ( x6 ) ;
assign n2638 =  ( n2615 ) ? ( n1071 ) : ( x6 ) ;
assign n2639 =  ( n2615 ) ? ( n1097 ) : ( x6 ) ;
assign n2640 =  ( n2615 ) ? ( n1105 ) : ( x6 ) ;
assign n2641 =  ( n2615 ) ? ( n1114 ) : ( x6 ) ;
assign n2642 =  ( n2615 ) ? ( n1120 ) : ( x6 ) ;
assign n2643 =  ( n2615 ) ? ( n1122 ) : ( x6 ) ;
assign n2644 =  ( n967 ) ? ( n2643 ) : ( x6 ) ;
assign n2645 =  ( n966 ) ? ( n2642 ) : ( n2644 ) ;
assign n2646 =  ( n965 ) ? ( n2641 ) : ( n2645 ) ;
assign n2647 =  ( n964 ) ? ( n2640 ) : ( n2646 ) ;
assign n2648 =  ( n963 ) ? ( n2639 ) : ( n2647 ) ;
assign n2649 =  ( n957 ) ? ( n2638 ) : ( n2648 ) ;
assign n2650 =  ( n956 ) ? ( n2637 ) : ( n2649 ) ;
assign n2651 =  ( n1068 ) ? ( n2636 ) : ( n2650 ) ;
assign n2652 =  ( n955 ) ? ( n2635 ) : ( n2651 ) ;
assign n2653 =  ( n954 ) ? ( n2633 ) : ( n2652 ) ;
assign n2654 =  ( n953 ) ? ( n2632 ) : ( n2653 ) ;
assign n2655 =  ( n952 ) ? ( n2631 ) : ( n2654 ) ;
assign n2656 =  ( n951 ) ? ( n2630 ) : ( n2655 ) ;
assign n2657 =  ( n950 ) ? ( n2629 ) : ( n2656 ) ;
assign n2658 =  ( n949 ) ? ( n2628 ) : ( n2657 ) ;
assign n2659 =  ( n947 ) ? ( n2627 ) : ( n2658 ) ;
assign n2660 =  ( n946 ) ? ( n2626 ) : ( n2659 ) ;
assign n2661 =  ( n943 ) ? ( n2625 ) : ( n2660 ) ;
assign n2662 =  ( n942 ) ? ( n2624 ) : ( n2661 ) ;
assign n2663 =  ( n939 ) ? ( n2623 ) : ( n2662 ) ;
assign n2664 =  ( n936 ) ? ( n2622 ) : ( n2663 ) ;
assign n2665 =  ( n934 ) ? ( n2621 ) : ( n2664 ) ;
assign n2666 =  ( n932 ) ? ( n2620 ) : ( n2665 ) ;
assign n2667 =  ( n930 ) ? ( n2619 ) : ( n2666 ) ;
assign n2668 =  ( n928 ) ? ( n2618 ) : ( n2667 ) ;
assign n2669 =  ( n926 ) ? ( n2617 ) : ( n2668 ) ;
assign n2670 =  ( n924 ) ? ( n2616 ) : ( n2669 ) ;
assign n2671 =  ( n621 ) ? ( n2670 ) : ( x6 ) ;
assign n2672 =  ( n1021 ) == ( 5'd7 )  ;
assign n2673 =  ( n2672 ) ? ( n1025 ) : ( x7 ) ;
assign n2674 =  ( n2672 ) ? ( n1027 ) : ( x7 ) ;
assign n2675 =  ( n2672 ) ? ( n1029 ) : ( x7 ) ;
assign n2676 =  ( n2672 ) ? ( n1031 ) : ( x7 ) ;
assign n2677 =  ( n2672 ) ? ( n1033 ) : ( x7 ) ;
assign n2678 =  ( n2672 ) ? ( n1035 ) : ( x7 ) ;
assign n2679 =  ( n2672 ) ? ( n1037 ) : ( x7 ) ;
assign n2680 =  ( n2672 ) ? ( n1039 ) : ( x7 ) ;
assign n2681 =  ( n2672 ) ? ( n1041 ) : ( x7 ) ;
assign n2682 =  ( n2672 ) ? ( n1043 ) : ( x7 ) ;
assign n2683 =  ( n2672 ) ? ( n1046 ) : ( x7 ) ;
assign n2684 =  ( n2672 ) ? ( n1048 ) : ( x7 ) ;
assign n2685 =  ( n2672 ) ? ( n1050 ) : ( x7 ) ;
assign n2686 =  ( n2672 ) ? ( n1053 ) : ( x7 ) ;
assign n2687 =  ( n2672 ) ? ( n1167 ) : ( x7 ) ;
assign n2688 =  ( n2672 ) ? ( n1058 ) : ( x7 ) ;
assign n2689 =  ( n2672 ) ? ( n1283 ) : ( x7 ) ;
assign n2690 =  ( n2672 ) ? ( n1064 ) : ( x7 ) ;
assign n2691 =  ( n2672 ) ? ( n1066 ) : ( x7 ) ;
assign n2692 =  ( n2672 ) ? ( n899 ) : ( x7 ) ;
assign n2693 =  ( n2672 ) ? ( n1072 ) : ( x7 ) ;
assign n2694 =  ( n2672 ) ? ( n1071 ) : ( x7 ) ;
assign n2695 =  ( n2672 ) ? ( n1097 ) : ( x7 ) ;
assign n2696 =  ( n2672 ) ? ( n1105 ) : ( x7 ) ;
assign n2697 =  ( n2672 ) ? ( n1114 ) : ( x7 ) ;
assign n2698 =  ( n2672 ) ? ( n1120 ) : ( x7 ) ;
assign n2699 =  ( n2672 ) ? ( n1122 ) : ( x7 ) ;
assign n2700 =  ( n967 ) ? ( n2699 ) : ( x7 ) ;
assign n2701 =  ( n966 ) ? ( n2698 ) : ( n2700 ) ;
assign n2702 =  ( n965 ) ? ( n2697 ) : ( n2701 ) ;
assign n2703 =  ( n964 ) ? ( n2696 ) : ( n2702 ) ;
assign n2704 =  ( n963 ) ? ( n2695 ) : ( n2703 ) ;
assign n2705 =  ( n957 ) ? ( n2694 ) : ( n2704 ) ;
assign n2706 =  ( n956 ) ? ( n2693 ) : ( n2705 ) ;
assign n2707 =  ( n1068 ) ? ( n2692 ) : ( n2706 ) ;
assign n2708 =  ( n955 ) ? ( n2691 ) : ( n2707 ) ;
assign n2709 =  ( n954 ) ? ( n2690 ) : ( n2708 ) ;
assign n2710 =  ( n953 ) ? ( n2689 ) : ( n2709 ) ;
assign n2711 =  ( n952 ) ? ( n2688 ) : ( n2710 ) ;
assign n2712 =  ( n951 ) ? ( n2687 ) : ( n2711 ) ;
assign n2713 =  ( n950 ) ? ( n2686 ) : ( n2712 ) ;
assign n2714 =  ( n949 ) ? ( n2685 ) : ( n2713 ) ;
assign n2715 =  ( n947 ) ? ( n2684 ) : ( n2714 ) ;
assign n2716 =  ( n946 ) ? ( n2683 ) : ( n2715 ) ;
assign n2717 =  ( n943 ) ? ( n2682 ) : ( n2716 ) ;
assign n2718 =  ( n942 ) ? ( n2681 ) : ( n2717 ) ;
assign n2719 =  ( n939 ) ? ( n2680 ) : ( n2718 ) ;
assign n2720 =  ( n936 ) ? ( n2679 ) : ( n2719 ) ;
assign n2721 =  ( n934 ) ? ( n2678 ) : ( n2720 ) ;
assign n2722 =  ( n932 ) ? ( n2677 ) : ( n2721 ) ;
assign n2723 =  ( n930 ) ? ( n2676 ) : ( n2722 ) ;
assign n2724 =  ( n928 ) ? ( n2675 ) : ( n2723 ) ;
assign n2725 =  ( n926 ) ? ( n2674 ) : ( n2724 ) ;
assign n2726 =  ( n924 ) ? ( n2673 ) : ( n2725 ) ;
assign n2727 =  ( n621 ) ? ( n2726 ) : ( x7 ) ;
assign n2728 =  ( n1021 ) == ( 5'd8 )  ;
assign n2729 =  ( n2728 ) ? ( n1025 ) : ( x8 ) ;
assign n2730 =  ( n2728 ) ? ( n1027 ) : ( x8 ) ;
assign n2731 =  ( n2728 ) ? ( n1029 ) : ( x8 ) ;
assign n2732 =  ( n2728 ) ? ( n1031 ) : ( x8 ) ;
assign n2733 =  ( n2728 ) ? ( n1033 ) : ( x8 ) ;
assign n2734 =  ( n2728 ) ? ( n1035 ) : ( x8 ) ;
assign n2735 =  ( n2728 ) ? ( n1037 ) : ( x8 ) ;
assign n2736 =  ( n2728 ) ? ( n1039 ) : ( x8 ) ;
assign n2737 =  ( n2728 ) ? ( n1041 ) : ( x8 ) ;
assign n2738 =  ( n2728 ) ? ( n1043 ) : ( x8 ) ;
assign n2739 =  ( n2728 ) ? ( n1046 ) : ( x8 ) ;
assign n2740 =  ( n2728 ) ? ( n1048 ) : ( x8 ) ;
assign n2741 =  ( n2728 ) ? ( n1050 ) : ( x8 ) ;
assign n2742 =  ( n2728 ) ? ( n1053 ) : ( x8 ) ;
assign n2743 =  ( n2728 ) ? ( n1167 ) : ( x8 ) ;
assign n2744 =  ( n2728 ) ? ( n1058 ) : ( x8 ) ;
assign n2745 =  ( n2728 ) ? ( n1283 ) : ( x8 ) ;
assign n2746 =  ( n2728 ) ? ( n1343 ) : ( x8 ) ;
assign n2747 =  ( n2728 ) ? ( n1066 ) : ( x8 ) ;
assign n2748 =  ( n2728 ) ? ( n899 ) : ( x8 ) ;
assign n2749 =  ( n2728 ) ? ( n1072 ) : ( x8 ) ;
assign n2750 =  ( n2728 ) ? ( n1071 ) : ( x8 ) ;
assign n2751 =  ( n2728 ) ? ( n1097 ) : ( x8 ) ;
assign n2752 =  ( n2728 ) ? ( n1105 ) : ( x8 ) ;
assign n2753 =  ( n2728 ) ? ( n1114 ) : ( x8 ) ;
assign n2754 =  ( n2728 ) ? ( n1120 ) : ( x8 ) ;
assign n2755 =  ( n2728 ) ? ( n1122 ) : ( x8 ) ;
assign n2756 =  ( n967 ) ? ( n2755 ) : ( x8 ) ;
assign n2757 =  ( n966 ) ? ( n2754 ) : ( n2756 ) ;
assign n2758 =  ( n965 ) ? ( n2753 ) : ( n2757 ) ;
assign n2759 =  ( n964 ) ? ( n2752 ) : ( n2758 ) ;
assign n2760 =  ( n963 ) ? ( n2751 ) : ( n2759 ) ;
assign n2761 =  ( n957 ) ? ( n2750 ) : ( n2760 ) ;
assign n2762 =  ( n956 ) ? ( n2749 ) : ( n2761 ) ;
assign n2763 =  ( n1068 ) ? ( n2748 ) : ( n2762 ) ;
assign n2764 =  ( n955 ) ? ( n2747 ) : ( n2763 ) ;
assign n2765 =  ( n954 ) ? ( n2746 ) : ( n2764 ) ;
assign n2766 =  ( n953 ) ? ( n2745 ) : ( n2765 ) ;
assign n2767 =  ( n952 ) ? ( n2744 ) : ( n2766 ) ;
assign n2768 =  ( n951 ) ? ( n2743 ) : ( n2767 ) ;
assign n2769 =  ( n950 ) ? ( n2742 ) : ( n2768 ) ;
assign n2770 =  ( n949 ) ? ( n2741 ) : ( n2769 ) ;
assign n2771 =  ( n947 ) ? ( n2740 ) : ( n2770 ) ;
assign n2772 =  ( n946 ) ? ( n2739 ) : ( n2771 ) ;
assign n2773 =  ( n943 ) ? ( n2738 ) : ( n2772 ) ;
assign n2774 =  ( n942 ) ? ( n2737 ) : ( n2773 ) ;
assign n2775 =  ( n939 ) ? ( n2736 ) : ( n2774 ) ;
assign n2776 =  ( n936 ) ? ( n2735 ) : ( n2775 ) ;
assign n2777 =  ( n934 ) ? ( n2734 ) : ( n2776 ) ;
assign n2778 =  ( n932 ) ? ( n2733 ) : ( n2777 ) ;
assign n2779 =  ( n930 ) ? ( n2732 ) : ( n2778 ) ;
assign n2780 =  ( n928 ) ? ( n2731 ) : ( n2779 ) ;
assign n2781 =  ( n926 ) ? ( n2730 ) : ( n2780 ) ;
assign n2782 =  ( n924 ) ? ( n2729 ) : ( n2781 ) ;
assign n2783 =  ( n621 ) ? ( n2782 ) : ( x8 ) ;
assign n2784 =  ( n1021 ) == ( 5'd9 )  ;
assign n2785 =  ( n2784 ) ? ( n1025 ) : ( x9 ) ;
assign n2786 =  ( n2784 ) ? ( n1027 ) : ( x9 ) ;
assign n2787 =  ( n2784 ) ? ( n1029 ) : ( x9 ) ;
assign n2788 =  ( n2784 ) ? ( n1031 ) : ( x9 ) ;
assign n2789 =  ( n2784 ) ? ( n1033 ) : ( x9 ) ;
assign n2790 =  ( n2784 ) ? ( n1035 ) : ( x9 ) ;
assign n2791 =  ( n2784 ) ? ( n1037 ) : ( x9 ) ;
assign n2792 =  ( n2784 ) ? ( n1039 ) : ( x9 ) ;
assign n2793 =  ( n2784 ) ? ( n1041 ) : ( x9 ) ;
assign n2794 =  ( n2784 ) ? ( n1043 ) : ( x9 ) ;
assign n2795 =  ( n2784 ) ? ( n1046 ) : ( x9 ) ;
assign n2796 =  ( n2784 ) ? ( n1048 ) : ( x9 ) ;
assign n2797 =  ( n2784 ) ? ( n1050 ) : ( x9 ) ;
assign n2798 =  ( n2784 ) ? ( n1452 ) : ( x9 ) ;
assign n2799 =  ( n2784 ) ? ( n1167 ) : ( x9 ) ;
assign n2800 =  ( n2784 ) ? ( n1058 ) : ( x9 ) ;
assign n2801 =  ( n2784 ) ? ( n1283 ) : ( x9 ) ;
assign n2802 =  ( n2784 ) ? ( n1343 ) : ( x9 ) ;
assign n2803 =  ( n2784 ) ? ( n1066 ) : ( x9 ) ;
assign n2804 =  ( n2784 ) ? ( n899 ) : ( x9 ) ;
assign n2805 =  ( n2784 ) ? ( n1072 ) : ( x9 ) ;
assign n2806 =  ( n2784 ) ? ( n1071 ) : ( x9 ) ;
assign n2807 =  ( n2784 ) ? ( n1097 ) : ( x9 ) ;
assign n2808 =  ( n2784 ) ? ( n1105 ) : ( x9 ) ;
assign n2809 =  ( n2784 ) ? ( n1114 ) : ( x9 ) ;
assign n2810 =  ( n2784 ) ? ( n1120 ) : ( x9 ) ;
assign n2811 =  ( n2784 ) ? ( n1122 ) : ( x9 ) ;
assign n2812 =  ( n967 ) ? ( n2811 ) : ( x9 ) ;
assign n2813 =  ( n966 ) ? ( n2810 ) : ( n2812 ) ;
assign n2814 =  ( n965 ) ? ( n2809 ) : ( n2813 ) ;
assign n2815 =  ( n964 ) ? ( n2808 ) : ( n2814 ) ;
assign n2816 =  ( n963 ) ? ( n2807 ) : ( n2815 ) ;
assign n2817 =  ( n957 ) ? ( n2806 ) : ( n2816 ) ;
assign n2818 =  ( n956 ) ? ( n2805 ) : ( n2817 ) ;
assign n2819 =  ( n1068 ) ? ( n2804 ) : ( n2818 ) ;
assign n2820 =  ( n955 ) ? ( n2803 ) : ( n2819 ) ;
assign n2821 =  ( n954 ) ? ( n2802 ) : ( n2820 ) ;
assign n2822 =  ( n953 ) ? ( n2801 ) : ( n2821 ) ;
assign n2823 =  ( n952 ) ? ( n2800 ) : ( n2822 ) ;
assign n2824 =  ( n951 ) ? ( n2799 ) : ( n2823 ) ;
assign n2825 =  ( n950 ) ? ( n2798 ) : ( n2824 ) ;
assign n2826 =  ( n949 ) ? ( n2797 ) : ( n2825 ) ;
assign n2827 =  ( n947 ) ? ( n2796 ) : ( n2826 ) ;
assign n2828 =  ( n946 ) ? ( n2795 ) : ( n2827 ) ;
assign n2829 =  ( n943 ) ? ( n2794 ) : ( n2828 ) ;
assign n2830 =  ( n942 ) ? ( n2793 ) : ( n2829 ) ;
assign n2831 =  ( n939 ) ? ( n2792 ) : ( n2830 ) ;
assign n2832 =  ( n936 ) ? ( n2791 ) : ( n2831 ) ;
assign n2833 =  ( n934 ) ? ( n2790 ) : ( n2832 ) ;
assign n2834 =  ( n932 ) ? ( n2789 ) : ( n2833 ) ;
assign n2835 =  ( n930 ) ? ( n2788 ) : ( n2834 ) ;
assign n2836 =  ( n928 ) ? ( n2787 ) : ( n2835 ) ;
assign n2837 =  ( n926 ) ? ( n2786 ) : ( n2836 ) ;
assign n2838 =  ( n924 ) ? ( n2785 ) : ( n2837 ) ;
assign n2839 =  ( n621 ) ? ( n2838 ) : ( x9 ) ;
assign n2840 =  ( 1'b1 ) & ( n620__take_int_or_expt )  ;
assign n2841 =  ( 1'b1 ) & ( n621 )  ;
assign n2842 = ~ ( n959 ) ;
assign n2843 =  ( n2841 ) & ( n2842 )  ;
assign n2844 = ~ ( n960 ) ;
assign n2845 =  ( n2843 ) & ( n2844 )  ;
assign n2846 = ~ ( n961 ) ;
assign n2847 =  ( n2845 ) & ( n2846 )  ;
assign n2848 =  ( n2845 ) & ( n961 )  ;
assign n2849 =  { ( n922 ) , ( n1021 ) }  ;
assign n2850 =  { {20{n2849[11] }  }, n2849}  ;
assign n2851 =  ( n807 ) + ( n2850 )  ;
assign n2852 = n2851[31:2] ;
assign n2853 =  {2'd0 , n2852}  ;
assign n2854 =  ( n888 ) & ( 32'd255 )  ;
assign n2855 = n2851[1:0] ;
assign n2856 =  {30'd0 , n2855}  ;
assign n2857 =  ( ( 32'd8 ) * ( n2856 ))  ;
assign n2858 =  ( n2854 ) << ( n2857 )  ;
assign n2859 =  ( 32'd255 ) << ( n2857 )  ;
assign n2860 = ~ ( n2859 ) ;
assign mem_addr_n2861 = n2853 ;
assign n2863 = mem_data_n2862 ;
assign n2864 =  ( n2860 ) & ( n2863 )  ;
assign n2865 =  ( n2858 ) | ( n2864 )  ;
assign n2866 =  ( n2843 ) & ( n960 )  ;
assign n2867 =  ( n888 ) & ( 32'd65535 )  ;
assign n2868 =  ( n2867 ) << ( n2857 )  ;
assign n2869 =  ( 32'd65535 ) << ( n2857 )  ;
assign n2870 = ~ ( n2869 ) ;
assign n2871 =  ( n2870 ) & ( n2863 )  ;
assign n2872 =  ( n2868 ) | ( n2871 )  ;
assign n2873 =  ( n2841 ) & ( n959 )  ;
assign n2874 =  ( n888 ) & ( 32'd4294967295 )  ;
assign n2875 =  ( n2874 ) << ( n2857 )  ;
assign n2876 =  ( 32'd4294967295 ) << ( n2857 )  ;
assign n2877 = ~ ( n2876 ) ;
assign n2878 =  ( n2877 ) & ( n2863 )  ;
assign n2879 =  ( n2875 ) | ( n2878 )  ;
assign mem_addr0 = n2873 ? (n2853) : (n2866 ? (n2853) : (n2848 ? (n2853) : (0)));
assign mem_data0 = n2873 ? (n2879) : (n2866 ? (n2872) : (n2848 ? (n2865) : ('dx)));
assign mem_wen0 = n2873 ? ( 1'b1 ) : (n2866 ? ( 1'b1 ) : (n2848 ? ( 1'b1 ) : (1'b0)));
always @(posedge clk) begin
   if(rst) begin
       Priv <= 2'd3;
       mbadaddr <= mbadaddr;
       mcause <= mcause;
       medeleg <= 32'd0;
       mepc <= mepc;
       mideleg <= 32'd0;
       mie <= 32'd0;
       mip <= 32'd0;
       misa <= 32'd1075052800;
       mscratch <= mscratch;
       mstatus <= 32'd0;
       mtvec <= 32'd0;
       pc <= pc;
       sbadaddr <= sbadaddr;
       scause <= scause;
       sepc <= sepc;
       sptbr <= 32'd0;
       sscratch <= sscratch;
       stvec <= 32'd0;
       x0 <= 32'd0;
       x1 <= x1;
       x10 <= x10;
       x11 <= x11;
       x12 <= x12;
       x13 <= x13;
       x14 <= x14;
       x15 <= x15;
       x16 <= x16;
       x17 <= x17;
       x18 <= x18;
       x19 <= x19;
       x2 <= x2;
       x20 <= x20;
       x21 <= x21;
       x22 <= x22;
       x23 <= x23;
       x24 <= x24;
       x25 <= x25;
       x26 <= x26;
       x27 <= x27;
       x28 <= x28;
       x29 <= x29;
       x3 <= x3;
       x30 <= x30;
       x31 <= x31;
       x4 <= x4;
       x5 <= x5;
       x6 <= x6;
       x7 <= x7;
       x8 <= x8;
       x9 <= x9;
   end
   else if(step) begin
       Priv <= n591;
       mbadaddr <= n623;
       mcause <= n671;
       medeleg <= n672;
       mepc <= n675;
       mideleg <= n676;
       mie <= n677;
       mip <= n17;
       misa <= n678;
       mscratch <= n679;
       mstatus <= n737;
       mtvec <= n738;
       pc <= n1007;
       sbadaddr <= n1010;
       scause <= n1015;
       sepc <= n1017;
       sptbr <= n1018;
       sscratch <= n1019;
       stvec <= n1020;
       x0 <= 32'd0;
       x1 <= n1151;
       x10 <= n1208;
       x11 <= n1264;
       x12 <= n1322;
       x13 <= n1381;
       x14 <= n1437;
       x15 <= n1494;
       x16 <= n1550;
       x17 <= n1606;
       x18 <= n1662;
       x19 <= n1718;
       x2 <= n1774;
       x20 <= n1830;
       x21 <= n1886;
       x22 <= n1942;
       x23 <= n1998;
       x24 <= n2054;
       x25 <= n2110;
       x26 <= n2166;
       x27 <= n2222;
       x28 <= n2278;
       x29 <= n2334;
       x3 <= n2390;
       x30 <= n2446;
       x31 <= n2502;
       x4 <= n2558;
       x5 <= n2614;
       x6 <= n2671;
       x7 <= n2727;
       x8 <= n2783;
       x9 <= n2839;
   end
end
endmodule
