module GB(
arg_0_TREADY,
arg_1_TDATA,
arg_1_TVALID,
LB1D_buff,
LB1D_in,
LB1D_it_1,
LB1D_p_cnt,
LB1D_uIn,
LB2D_proc_w,
LB2D_proc_x,
LB2D_proc_y,
LB2D_shift_0,
LB2D_shift_1,
LB2D_shift_2,
LB2D_shift_3,
LB2D_shift_4,
LB2D_shift_5,
LB2D_shift_6,
LB2D_shift_7,
LB2D_shift_x,
LB2D_shift_y,
arg_0_TDATA,
arg_0_TVALID,
arg_1_TREADY,
gb_exit_it_1,
gb_exit_it_2,
gb_exit_it_3,
gb_exit_it_4,
gb_exit_it_5,
gb_exit_it_6,
gb_exit_it_7,
gb_exit_it_8,
gb_p_cnt,
gb_pp_it_1,
gb_pp_it_2,
gb_pp_it_3,
gb_pp_it_4,
gb_pp_it_5,
gb_pp_it_6,
gb_pp_it_7,
gb_pp_it_8,
gb_pp_it_9,
in_stream_buff_0,
in_stream_buff_1,
in_stream_empty,
in_stream_full,
slice_stream_buff_0,
slice_stream_buff_1,
slice_stream_empty,
slice_stream_full,
stencil_stream_buff_0,
stencil_stream_buff_1,
stencil_stream_empty,
stencil_stream_full,
clk,rst,
step
);
input            arg_0_TREADY;
input      [7:0] arg_1_TDATA;
input            arg_1_TVALID;
input clk;
input rst;
input step;
output      [7:0] LB1D_buff;
output      [7:0] LB1D_in;
output            LB1D_it_1;
output     [18:0] LB1D_p_cnt;
output      [7:0] LB1D_uIn;
output     [63:0] LB2D_proc_w;
output      [8:0] LB2D_proc_x;
output      [9:0] LB2D_proc_y;
output     [71:0] LB2D_shift_0;
output     [71:0] LB2D_shift_1;
output     [71:0] LB2D_shift_2;
output     [71:0] LB2D_shift_3;
output     [71:0] LB2D_shift_4;
output     [71:0] LB2D_shift_5;
output     [71:0] LB2D_shift_6;
output     [71:0] LB2D_shift_7;
output      [8:0] LB2D_shift_x;
output      [9:0] LB2D_shift_y;
output      [7:0] arg_0_TDATA;
output            arg_0_TVALID;
output            arg_1_TREADY;
output            gb_exit_it_1;
output            gb_exit_it_2;
output            gb_exit_it_3;
output            gb_exit_it_4;
output            gb_exit_it_5;
output            gb_exit_it_6;
output            gb_exit_it_7;
output            gb_exit_it_8;
output     [18:0] gb_p_cnt;
output            gb_pp_it_1;
output            gb_pp_it_2;
output            gb_pp_it_3;
output            gb_pp_it_4;
output            gb_pp_it_5;
output            gb_pp_it_6;
output            gb_pp_it_7;
output            gb_pp_it_8;
output            gb_pp_it_9;
output      [7:0] in_stream_buff_0;
output      [7:0] in_stream_buff_1;
output            in_stream_empty;
output            in_stream_full;
output     [71:0] slice_stream_buff_0;
output     [71:0] slice_stream_buff_1;
output            slice_stream_empty;
output            slice_stream_full;
output    [647:0] stencil_stream_buff_0;
output    [647:0] stencil_stream_buff_1;
output            stencil_stream_empty;
output            stencil_stream_full;
reg      [7:0] LB1D_buff;
reg      [7:0] LB1D_in;
reg            LB1D_it_1;
reg     [18:0] LB1D_p_cnt;
reg      [7:0] LB1D_uIn;
reg     [63:0] LB2D_proc_w;
reg      [8:0] LB2D_proc_x;
reg      [9:0] LB2D_proc_y;
reg     [71:0] LB2D_shift_0;
reg     [71:0] LB2D_shift_1;
reg     [71:0] LB2D_shift_2;
reg     [71:0] LB2D_shift_3;
reg     [71:0] LB2D_shift_4;
reg     [71:0] LB2D_shift_5;
reg     [71:0] LB2D_shift_6;
reg     [71:0] LB2D_shift_7;
reg      [8:0] LB2D_shift_x;
reg      [9:0] LB2D_shift_y;
reg      [7:0] arg_0_TDATA;
reg            arg_0_TVALID;
reg            arg_1_TREADY;
reg            gb_exit_it_1;
reg            gb_exit_it_2;
reg            gb_exit_it_3;
reg            gb_exit_it_4;
reg            gb_exit_it_5;
reg            gb_exit_it_6;
reg            gb_exit_it_7;
reg            gb_exit_it_8;
reg     [18:0] gb_p_cnt;
reg            gb_pp_it_1;
reg            gb_pp_it_2;
reg            gb_pp_it_3;
reg            gb_pp_it_4;
reg            gb_pp_it_5;
reg            gb_pp_it_6;
reg            gb_pp_it_7;
reg            gb_pp_it_8;
reg            gb_pp_it_9;
reg      [7:0] in_stream_buff_0;
reg      [7:0] in_stream_buff_1;
reg            in_stream_empty;
reg            in_stream_full;
reg     [71:0] slice_stream_buff_0;
reg     [71:0] slice_stream_buff_1;
reg            slice_stream_empty;
reg            slice_stream_full;
reg    [647:0] stencil_stream_buff_0;
reg    [647:0] stencil_stream_buff_1;
reg            stencil_stream_empty;
reg            stencil_stream_full;
wire            arg_0_TREADY;
wire      [7:0] arg_1_TDATA;
wire            arg_1_TVALID;
wire            n0;
wire            n1;
wire            n2;
wire            n3;
wire            n4;
wire            n5;
wire            n6;
wire            n7;
wire            n8;
wire            n9;
wire            n10;
wire            n11;
wire            n12;
wire            n13;
wire            n14;
wire            n15;
wire            n16;
wire            n17;
wire            n18;
wire            n19;
wire            n20;
wire            n21;
wire            n22;
wire            n23;
wire            n24;
wire            n25;
wire            n26;
wire            n27;
wire            n28;
wire            n29;
wire            n30;
wire            n31;
wire            n32;
wire            n33;
wire            n34;
wire            n35;
wire            n36;
wire            n37;
wire      [7:0] n38;
wire      [7:0] n39;
wire      [7:0] n40;
wire      [7:0] n41;
wire      [7:0] n42;
wire      [7:0] n43;
wire      [7:0] n44;
wire      [7:0] n45;
wire      [7:0] n46;
wire      [7:0] n47;
wire      [7:0] n48;
wire      [7:0] n49;
wire            n50;
wire            n51;
wire            n52;
wire     [18:0] n53;
wire     [18:0] n54;
wire            n55;
wire     [18:0] n56;
wire     [18:0] n57;
wire     [18:0] n58;
wire     [18:0] n59;
wire     [18:0] n60;
wire     [18:0] n61;
wire     [18:0] n62;
wire     [18:0] n63;
wire      [7:0] n64;
wire      [7:0] n65;
wire      [7:0] n66;
wire      [7:0] n67;
wire      [7:0] n68;
wire            n69;
wire            n70;
wire            n71;
wire            n72;
wire     [63:0] n73;
wire     [63:0] n74;
wire     [63:0] n75;
wire     [63:0] n76;
wire     [63:0] n77;
wire     [63:0] n78;
wire     [63:0] n79;
wire     [63:0] n80;
wire     [63:0] n81;
wire            n82;
wire      [8:0] n83;
wire      [8:0] n84;
wire      [8:0] n85;
wire      [8:0] n86;
wire      [8:0] n87;
wire      [8:0] n88;
wire      [8:0] n89;
wire      [8:0] n90;
wire      [8:0] n91;
wire            n92;
wire      [9:0] n93;
wire      [9:0] n94;
wire      [9:0] n95;
wire      [9:0] n96;
wire      [9:0] n97;
wire      [9:0] n98;
wire      [9:0] n99;
wire      [9:0] n100;
wire      [9:0] n101;
wire            n102;
wire     [71:0] n103;
wire     [71:0] n104;
wire     [71:0] n105;
wire     [71:0] n106;
wire     [71:0] n107;
wire     [71:0] n108;
wire     [71:0] n109;
wire     [71:0] n110;
wire     [71:0] n111;
wire     [71:0] n112;
wire     [71:0] n113;
wire     [71:0] n114;
wire     [71:0] n115;
wire     [71:0] n116;
wire     [71:0] n117;
wire     [71:0] n118;
wire     [71:0] n119;
wire     [71:0] n120;
wire     [71:0] n121;
wire     [71:0] n122;
wire     [71:0] n123;
wire     [71:0] n124;
wire     [71:0] n125;
wire     [71:0] n126;
wire     [71:0] n127;
wire     [71:0] n128;
wire     [71:0] n129;
wire     [71:0] n130;
wire     [71:0] n131;
wire     [71:0] n132;
wire     [71:0] n133;
wire     [71:0] n134;
wire     [71:0] n135;
wire     [71:0] n136;
wire     [71:0] n137;
wire     [71:0] n138;
wire     [71:0] n139;
wire     [71:0] n140;
wire     [71:0] n141;
wire     [71:0] n142;
wire     [71:0] n143;
wire     [71:0] n144;
wire     [71:0] n145;
wire     [71:0] n146;
wire     [71:0] n147;
wire     [71:0] n148;
wire     [71:0] n149;
wire     [71:0] n150;
wire     [71:0] n151;
wire      [8:0] n152;
wire      [8:0] n153;
wire      [8:0] n154;
wire      [8:0] n155;
wire      [8:0] n156;
wire      [8:0] n157;
wire      [8:0] n158;
wire            n159;
wire            n160;
wire      [9:0] n161;
wire      [9:0] n162;
wire      [9:0] n163;
wire      [9:0] n164;
wire      [9:0] n165;
wire      [9:0] n166;
wire      [9:0] n167;
wire      [9:0] n168;
wire      [9:0] n169;
wire            n170;
wire    [647:0] n171;
wire      [7:0] n172;
wire      [7:0] n173;
wire      [7:0] n174;
wire      [7:0] n175;
wire      [7:0] n176;
wire      [7:0] n177;
wire      [7:0] n178;
wire            n179;
wire            n180;
wire            n181;
wire            n182;
wire            n183;
wire            n184;
wire            n185;
wire            n186;
wire            n187;
wire            n188;
wire            n189;
wire            n190;
wire            n191;
wire            n192;
wire            n193;
wire     [18:0] n194;
wire            n195;
wire            n196;
wire            n197;
wire            n198;
wire            n199;
wire            n200;
wire            n201;
wire            n202;
wire            n203;
wire            n204;
wire            n205;
wire            n206;
wire            n207;
wire            n208;
wire            n209;
wire            n210;
wire            n211;
wire            n212;
wire            n213;
wire            n214;
wire            n215;
wire            n216;
wire            n217;
wire            n218;
wire            n219;
wire            n220;
wire            n221;
wire            n222;
wire            n223;
wire            n224;
wire            n225;
wire            n226;
wire            n227;
wire            n228;
wire            n229;
wire            n230;
wire            n231;
wire            n232;
wire            n233;
wire            n234;
wire            n235;
wire            n236;
wire            n237;
wire            n238;
wire            n239;
wire            n240;
wire            n241;
wire            n242;
wire            n243;
wire            n244;
wire            n245;
wire     [18:0] n246;
wire     [18:0] n247;
wire     [18:0] n248;
wire     [18:0] n249;
wire     [18:0] n250;
wire     [18:0] n251;
wire     [18:0] n252;
wire            n253;
wire            n254;
wire            n255;
wire            n256;
wire            n257;
wire            n258;
wire            n259;
wire            n260;
wire            n261;
wire            n262;
wire            n263;
wire            n264;
wire            n265;
wire            n266;
wire            n267;
wire            n268;
wire            n269;
wire            n270;
wire            n271;
wire            n272;
wire            n273;
wire            n274;
wire            n275;
wire            n276;
wire            n277;
wire            n278;
wire            n279;
wire            n280;
wire            n281;
wire            n282;
wire            n283;
wire            n284;
wire            n285;
wire            n286;
wire            n287;
wire            n288;
wire            n289;
wire            n290;
wire            n291;
wire            n292;
wire            n293;
wire            n294;
wire            n295;
wire            n296;
wire            n297;
wire            n298;
wire            n299;
wire            n300;
wire            n301;
wire            n302;
wire            n303;
wire            n304;
wire            n305;
wire            n306;
wire      [7:0] n307;
wire      [7:0] n308;
wire      [7:0] n309;
wire      [7:0] n310;
wire      [7:0] n311;
wire      [7:0] n312;
wire      [7:0] n313;
wire      [7:0] n314;
wire      [7:0] n315;
wire      [7:0] n316;
wire      [7:0] n317;
wire      [7:0] n318;
wire            n319;
wire            n320;
wire            n321;
wire            n322;
wire            n323;
wire            n324;
wire            n325;
wire            n326;
wire            n327;
wire            n328;
wire            n329;
wire            n330;
wire            n331;
wire            n332;
wire            n333;
wire            n334;
wire      [7:0] n335;
wire            n336;
wire      [7:0] n337;
wire            n338;
wire      [7:0] n339;
wire            n340;
wire      [7:0] n341;
wire            n342;
wire      [7:0] n343;
wire            n344;
wire      [7:0] n345;
wire            n346;
wire      [7:0] n347;
wire            n348;
wire      [7:0] n349;
wire      [7:0] n350;
wire      [7:0] n351;
wire      [7:0] n352;
wire      [7:0] n353;
wire      [7:0] n354;
wire      [7:0] n355;
wire      [7:0] n356;
wire      [7:0] n357;
wire      [7:0] n358;
wire      [7:0] n359;
wire      [7:0] n360;
wire      [7:0] n361;
wire      [7:0] n362;
wire      [7:0] n363;
wire      [7:0] n364;
wire      [7:0] n365;
wire      [7:0] n366;
wire      [7:0] n367;
wire      [7:0] n368;
wire      [7:0] n369;
wire      [7:0] n370;
wire      [7:0] n371;
wire      [7:0] n372;
wire      [7:0] n373;
wire      [7:0] n374;
wire      [7:0] n375;
wire      [7:0] n376;
wire      [7:0] n377;
wire      [7:0] n378;
wire      [7:0] n379;
wire      [7:0] n380;
wire      [7:0] n381;
wire      [7:0] n382;
wire      [7:0] n383;
wire      [7:0] n384;
wire      [7:0] n385;
wire      [7:0] n386;
wire      [7:0] n387;
wire      [7:0] n388;
wire      [7:0] n389;
wire      [7:0] n390;
wire      [7:0] n391;
wire      [7:0] n392;
wire      [7:0] n393;
wire      [7:0] n394;
wire      [7:0] n395;
wire      [7:0] n396;
wire      [7:0] n397;
wire      [7:0] n398;
wire      [7:0] n399;
wire      [7:0] n400;
wire      [7:0] n401;
wire      [7:0] n402;
wire      [7:0] n403;
wire      [7:0] n404;
wire      [7:0] n405;
wire      [7:0] n406;
wire     [15:0] n407;
wire     [23:0] n408;
wire     [31:0] n409;
wire     [39:0] n410;
wire     [47:0] n411;
wire     [55:0] n412;
wire     [63:0] n413;
wire     [71:0] n414;
wire     [71:0] n415;
wire     [71:0] n416;
wire     [71:0] n417;
wire     [71:0] n418;
wire     [71:0] n419;
wire     [71:0] n420;
wire     [71:0] n421;
wire     [71:0] n422;
wire     [71:0] n423;
wire     [71:0] n424;
wire     [71:0] n425;
wire     [71:0] n426;
wire     [71:0] n427;
wire     [71:0] n428;
wire            n429;
wire            n430;
wire            n431;
wire            n432;
wire            n433;
wire            n434;
wire            n435;
wire            n436;
wire            n437;
wire            n438;
wire            n439;
wire            n440;
wire            n441;
wire            n442;
wire            n443;
wire            n444;
wire            n445;
wire            n446;
wire      [7:0] n447;
wire      [7:0] n448;
wire      [7:0] n449;
wire      [7:0] n450;
wire      [7:0] n451;
wire      [7:0] n452;
wire      [7:0] n453;
wire      [7:0] n454;
wire      [7:0] n455;
wire     [15:0] n456;
wire     [23:0] n457;
wire     [31:0] n458;
wire     [39:0] n459;
wire     [47:0] n460;
wire     [55:0] n461;
wire     [63:0] n462;
wire     [71:0] n463;
wire      [7:0] n464;
wire      [7:0] n465;
wire      [7:0] n466;
wire      [7:0] n467;
wire      [7:0] n468;
wire      [7:0] n469;
wire      [7:0] n470;
wire      [7:0] n471;
wire      [7:0] n472;
wire     [15:0] n473;
wire     [23:0] n474;
wire     [31:0] n475;
wire     [39:0] n476;
wire     [47:0] n477;
wire     [55:0] n478;
wire     [63:0] n479;
wire     [71:0] n480;
wire      [7:0] n481;
wire      [7:0] n482;
wire      [7:0] n483;
wire      [7:0] n484;
wire      [7:0] n485;
wire      [7:0] n486;
wire      [7:0] n487;
wire      [7:0] n488;
wire      [7:0] n489;
wire     [15:0] n490;
wire     [23:0] n491;
wire     [31:0] n492;
wire     [39:0] n493;
wire     [47:0] n494;
wire     [55:0] n495;
wire     [63:0] n496;
wire     [71:0] n497;
wire      [7:0] n498;
wire      [7:0] n499;
wire      [7:0] n500;
wire      [7:0] n501;
wire      [7:0] n502;
wire      [7:0] n503;
wire      [7:0] n504;
wire      [7:0] n505;
wire      [7:0] n506;
wire     [15:0] n507;
wire     [23:0] n508;
wire     [31:0] n509;
wire     [39:0] n510;
wire     [47:0] n511;
wire     [55:0] n512;
wire     [63:0] n513;
wire     [71:0] n514;
wire      [7:0] n515;
wire      [7:0] n516;
wire      [7:0] n517;
wire      [7:0] n518;
wire      [7:0] n519;
wire      [7:0] n520;
wire      [7:0] n521;
wire      [7:0] n522;
wire      [7:0] n523;
wire     [15:0] n524;
wire     [23:0] n525;
wire     [31:0] n526;
wire     [39:0] n527;
wire     [47:0] n528;
wire     [55:0] n529;
wire     [63:0] n530;
wire     [71:0] n531;
wire      [7:0] n532;
wire      [7:0] n533;
wire      [7:0] n534;
wire      [7:0] n535;
wire      [7:0] n536;
wire      [7:0] n537;
wire      [7:0] n538;
wire      [7:0] n539;
wire      [7:0] n540;
wire     [15:0] n541;
wire     [23:0] n542;
wire     [31:0] n543;
wire     [39:0] n544;
wire     [47:0] n545;
wire     [55:0] n546;
wire     [63:0] n547;
wire     [71:0] n548;
wire      [7:0] n549;
wire      [7:0] n550;
wire      [7:0] n551;
wire      [7:0] n552;
wire      [7:0] n553;
wire      [7:0] n554;
wire      [7:0] n555;
wire      [7:0] n556;
wire      [7:0] n557;
wire     [15:0] n558;
wire     [23:0] n559;
wire     [31:0] n560;
wire     [39:0] n561;
wire     [47:0] n562;
wire     [55:0] n563;
wire     [63:0] n564;
wire     [71:0] n565;
wire      [7:0] n566;
wire      [7:0] n567;
wire      [7:0] n568;
wire      [7:0] n569;
wire      [7:0] n570;
wire      [7:0] n571;
wire      [7:0] n572;
wire      [7:0] n573;
wire      [7:0] n574;
wire     [15:0] n575;
wire     [23:0] n576;
wire     [31:0] n577;
wire     [39:0] n578;
wire     [47:0] n579;
wire     [55:0] n580;
wire     [63:0] n581;
wire     [71:0] n582;
wire      [7:0] n583;
wire      [7:0] n584;
wire      [7:0] n585;
wire      [7:0] n586;
wire      [7:0] n587;
wire      [7:0] n588;
wire      [7:0] n589;
wire      [7:0] n590;
wire      [7:0] n591;
wire     [15:0] n592;
wire     [23:0] n593;
wire     [31:0] n594;
wire     [39:0] n595;
wire     [47:0] n596;
wire     [55:0] n597;
wire     [63:0] n598;
wire     [71:0] n599;
wire    [143:0] n600;
wire    [215:0] n601;
wire    [287:0] n602;
wire    [359:0] n603;
wire    [431:0] n604;
wire    [503:0] n605;
wire    [575:0] n606;
wire    [647:0] n607;
wire    [647:0] n608;
wire    [647:0] n609;
wire    [647:0] n610;
wire    [647:0] n611;
wire    [647:0] n612;
wire    [647:0] n613;
wire    [647:0] n614;
wire    [647:0] n615;
wire    [647:0] n616;
wire    [647:0] n617;
wire    [647:0] n618;
wire    [647:0] n619;
wire    [647:0] n620;
wire            n621;
wire            n622;
wire            n623;
wire            n624;
wire            n625;
wire            n626;
wire            n627;
wire            n628;
wire            n629;
wire            n630;
wire            n631;
wire            n632;
wire            n633;
wire            n634;
wire            n635;
wire            n636;
wire            n637;
wire            n638;
wire      [8:0] LB2D_proc_0_addr0;
wire      [7:0] LB2D_proc_0_data0;
wire            n639;
wire            n640;
wire            n641;
wire            n642;
wire            n643;
wire            n644;
wire            n645;
wire            n646;
wire            n647;
wire            n648;
wire            n649;
wire            n650;
wire            n651;
wire            n652;
wire            n653;
wire            n654;
wire            n655;
wire            n656;
wire            n657;
wire      [8:0] LB2D_proc_1_addr0;
wire      [7:0] LB2D_proc_1_data0;
wire            n658;
wire            n659;
wire            n660;
wire      [8:0] LB2D_proc_2_addr0;
wire      [7:0] LB2D_proc_2_data0;
wire            n661;
wire            n662;
wire            n663;
wire      [8:0] LB2D_proc_3_addr0;
wire      [7:0] LB2D_proc_3_data0;
wire            n664;
wire            n665;
wire            n666;
wire      [8:0] LB2D_proc_4_addr0;
wire      [7:0] LB2D_proc_4_data0;
wire            n667;
wire            n668;
wire            n669;
wire      [8:0] LB2D_proc_5_addr0;
wire      [7:0] LB2D_proc_5_data0;
wire            n670;
wire            n671;
wire            n672;
wire      [8:0] LB2D_proc_6_addr0;
wire      [7:0] LB2D_proc_6_data0;
wire            n673;
wire            n674;
wire            n675;
wire      [8:0] LB2D_proc_7_addr0;
wire      [7:0] LB2D_proc_7_data0;
wire            n676;
wire            n677;
wire            n678;
reg      [7:0] LB2D_proc_0[511:0];
reg      [7:0] LB2D_proc_1[511:0];
reg      [7:0] LB2D_proc_2[511:0];
reg      [7:0] LB2D_proc_3[511:0];
reg      [7:0] LB2D_proc_4[511:0];
reg      [7:0] LB2D_proc_5[511:0];
reg      [7:0] LB2D_proc_6[511:0];
reg      [7:0] LB2D_proc_7[511:0];
wire clk;
wire rst;
wire step;
assign n0 =  ( arg_0_TREADY ) == ( 1'd1 )  ;
assign n1 =  ( arg_0_TVALID ) == ( 1'd1 )  ;
assign n2 =  ( n0 ) & ( n1 )  ;
assign n3 =  ( arg_1_TVALID ) == ( 1'd0 )  ;
assign n4 =  ( n2 ) & ( n3 )  ;
assign n5 =  ( arg_1_TREADY ) == ( 1'd1 )  ;
assign n6 =  ( arg_1_TVALID ) == ( 1'd1 )  ;
assign n7 =  ( n5 ) & ( n6 )  ;
assign n8 =  ( arg_0_TREADY ) == ( 1'd0 )  ;
assign n9 =  ( n7 ) & ( n8 )  ;
assign n10 =  ( arg_0_TVALID ) == ( 1'd0 )  ;
assign n11 =  ( gb_exit_it_1 ) == ( 1'd0 )  ;
assign n12 =  ( stencil_stream_empty ) == ( 1'd0 )  ;
assign n13 =  ( n11 ) & ( n12 )  ;
assign n14 =  ( gb_exit_it_1 ) == ( 1'd1 )  ;
assign n15 =  ( gb_exit_it_8 ) == ( 1'd0 )  ;
assign n16 =  ( n14 ) & ( n15 )  ;
assign n17 =  ( n13 ) | ( n16 )  ;
assign n18 =  ( n10 ) & ( n17 )  ;
assign n19 =  ( slice_stream_empty ) == ( 1'd0 )  ;
assign n20 =  ( LB2D_shift_x ) != ( 9'd488 )  ;
assign n21 =  ( n19 ) & ( n20 )  ;
assign n22 =  ( stencil_stream_full ) == ( 1'd0 )  ;
assign n23 =  ( LB2D_shift_x ) < ( 9'd8 )  ;
assign n24 =  ( n22 ) | ( n23 )  ;
assign n25 =  ( n21 ) & ( n24 )  ;
assign n26 =  ( in_stream_empty ) == ( 1'd0 )  ;
assign n27 =  ( LB2D_proc_x ) != ( 9'd488 )  ;
assign n28 =  ( n26 ) & ( n27 )  ;
assign n29 =  ( slice_stream_full ) == ( 1'd0 )  ;
assign n30 =  ( LB2D_proc_y ) < ( 10'd8 )  ;
assign n31 =  ( n29 ) | ( n30 )  ;
assign n32 =  ( n28 ) & ( n31 )  ;
assign n33 =  ( arg_1_TREADY ) == ( 1'd0 )  ;
assign n34 =  ( in_stream_full ) == ( 1'd0 )  ;
assign n35 =  ( n33 ) & ( n34 )  ;
assign n36 =  ( LB1D_it_1 ) == ( 1'd1 )  ;
assign n37 =  ( n35 ) & ( n36 )  ;
assign n38 =  ( n37 ) ? ( LB1D_uIn ) : ( LB1D_buff ) ;
assign n39 =  ( n32 ) ? ( LB1D_buff ) : ( n38 ) ;
assign n40 =  ( n25 ) ? ( LB1D_buff ) : ( n39 ) ;
assign n41 =  ( n18 ) ? ( LB1D_buff ) : ( n40 ) ;
assign n42 =  ( n9 ) ? ( LB1D_buff ) : ( n41 ) ;
assign n43 =  ( n4 ) ? ( LB1D_buff ) : ( n42 ) ;
assign n44 =  ( n37 ) ? ( LB1D_in ) : ( LB1D_in ) ;
assign n45 =  ( n32 ) ? ( LB1D_in ) : ( n44 ) ;
assign n46 =  ( n25 ) ? ( LB1D_in ) : ( n45 ) ;
assign n47 =  ( n18 ) ? ( LB1D_in ) : ( n46 ) ;
assign n48 =  ( n9 ) ? ( arg_1_TDATA ) : ( n47 ) ;
assign n49 =  ( n4 ) ? ( LB1D_in ) : ( n48 ) ;
assign n50 =  ( LB1D_it_1 ) == ( 1'd0 )  ;
assign n51 =  ( n35 ) & ( n50 )  ;
assign n52 =  ( n51 ) ? ( 1'd1 ) : ( LB1D_it_1 ) ;
assign n53 =  ( LB1D_p_cnt ) + ( 19'd1 )  ;
assign n54 =  ( 19'd316224 ) - ( 19'd1 )  ;
assign n55 =  ( LB1D_p_cnt ) == ( n54 )  ;
assign n56 =  ( n55 ) ? ( 19'd0 ) : ( n53 ) ;
assign n57 =  ( n37 ) ? ( n56 ) : ( LB1D_p_cnt ) ;
assign n58 =  ( n51 ) ? ( n53 ) : ( n57 ) ;
assign n59 =  ( n32 ) ? ( LB1D_p_cnt ) : ( n58 ) ;
assign n60 =  ( n25 ) ? ( LB1D_p_cnt ) : ( n59 ) ;
assign n61 =  ( n18 ) ? ( LB1D_p_cnt ) : ( n60 ) ;
assign n62 =  ( n9 ) ? ( LB1D_p_cnt ) : ( n61 ) ;
assign n63 =  ( n4 ) ? ( LB1D_p_cnt ) : ( n62 ) ;
assign n64 =  ( n37 ) ? ( LB1D_in ) : ( LB1D_uIn ) ;
assign n65 =  ( n32 ) ? ( LB1D_uIn ) : ( n64 ) ;
assign n66 =  ( n25 ) ? ( LB1D_uIn ) : ( n65 ) ;
assign n67 =  ( n18 ) ? ( LB1D_uIn ) : ( n66 ) ;
assign n68 =  ( n9 ) ? ( LB1D_uIn ) : ( n67 ) ;
assign n69 =  ( LB2D_proc_x ) == ( 9'd488 )  ;
assign n70 =  ( n26 ) & ( n69 )  ;
assign n71 =  ( n70 ) & ( n31 )  ;
assign n72 =  ( LB2D_proc_w ) == ( 64'd7 )  ;
assign n73 =  ( LB2D_proc_w ) + ( 64'd1 )  ;
assign n74 =  ( n72 ) ? ( 64'd0 ) : ( n73 ) ;
assign n75 =  ( n37 ) ? ( LB2D_proc_w ) : ( LB2D_proc_w ) ;
assign n76 =  ( n32 ) ? ( LB2D_proc_w ) : ( n75 ) ;
assign n77 =  ( n71 ) ? ( n74 ) : ( n76 ) ;
assign n78 =  ( n25 ) ? ( LB2D_proc_w ) : ( n77 ) ;
assign n79 =  ( n18 ) ? ( LB2D_proc_w ) : ( n78 ) ;
assign n80 =  ( n9 ) ? ( LB2D_proc_w ) : ( n79 ) ;
assign n81 =  ( n4 ) ? ( LB2D_proc_w ) : ( n80 ) ;
assign n82 =  ( LB2D_proc_x ) == ( 9'd0 )  ;
assign n83 =  ( LB2D_proc_x ) + ( 9'd1 )  ;
assign n84 =  ( n82 ) ? ( 9'd1 ) : ( n83 ) ;
assign n85 =  ( n37 ) ? ( LB2D_proc_x ) : ( LB2D_proc_x ) ;
assign n86 =  ( n32 ) ? ( n84 ) : ( n85 ) ;
assign n87 =  ( n71 ) ? ( 9'd0 ) : ( n86 ) ;
assign n88 =  ( n25 ) ? ( LB2D_proc_x ) : ( n87 ) ;
assign n89 =  ( n18 ) ? ( LB2D_proc_x ) : ( n88 ) ;
assign n90 =  ( n9 ) ? ( LB2D_proc_x ) : ( n89 ) ;
assign n91 =  ( n4 ) ? ( LB2D_proc_x ) : ( n90 ) ;
assign n92 =  ( LB2D_proc_y ) == ( 10'd488 )  ;
assign n93 =  ( LB2D_proc_y ) + ( 10'd1 )  ;
assign n94 =  ( n92 ) ? ( 10'd0 ) : ( n93 ) ;
assign n95 =  ( n37 ) ? ( LB2D_proc_y ) : ( LB2D_proc_y ) ;
assign n96 =  ( n32 ) ? ( LB2D_proc_y ) : ( n95 ) ;
assign n97 =  ( n71 ) ? ( n94 ) : ( n96 ) ;
assign n98 =  ( n25 ) ? ( LB2D_proc_y ) : ( n97 ) ;
assign n99 =  ( n18 ) ? ( LB2D_proc_y ) : ( n98 ) ;
assign n100 =  ( n9 ) ? ( LB2D_proc_y ) : ( n99 ) ;
assign n101 =  ( n4 ) ? ( LB2D_proc_y ) : ( n100 ) ;
assign n102 =  ( slice_stream_full ) == ( 1'd1 )  ;
assign n103 =  ( n102 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n104 =  ( n37 ) ? ( LB2D_shift_0 ) : ( LB2D_shift_0 ) ;
assign n105 =  ( n32 ) ? ( LB2D_shift_0 ) : ( n104 ) ;
assign n106 =  ( n25 ) ? ( n103 ) : ( n105 ) ;
assign n107 =  ( n18 ) ? ( LB2D_shift_0 ) : ( n106 ) ;
assign n108 =  ( n9 ) ? ( LB2D_shift_0 ) : ( n107 ) ;
assign n109 =  ( n4 ) ? ( LB2D_shift_0 ) : ( n108 ) ;
assign n110 =  ( n37 ) ? ( LB2D_shift_1 ) : ( LB2D_shift_1 ) ;
assign n111 =  ( n32 ) ? ( LB2D_shift_1 ) : ( n110 ) ;
assign n112 =  ( n25 ) ? ( LB2D_shift_0 ) : ( n111 ) ;
assign n113 =  ( n18 ) ? ( LB2D_shift_1 ) : ( n112 ) ;
assign n114 =  ( n9 ) ? ( LB2D_shift_1 ) : ( n113 ) ;
assign n115 =  ( n4 ) ? ( LB2D_shift_1 ) : ( n114 ) ;
assign n116 =  ( n37 ) ? ( LB2D_shift_2 ) : ( LB2D_shift_2 ) ;
assign n117 =  ( n32 ) ? ( LB2D_shift_2 ) : ( n116 ) ;
assign n118 =  ( n25 ) ? ( LB2D_shift_1 ) : ( n117 ) ;
assign n119 =  ( n18 ) ? ( LB2D_shift_2 ) : ( n118 ) ;
assign n120 =  ( n9 ) ? ( LB2D_shift_2 ) : ( n119 ) ;
assign n121 =  ( n4 ) ? ( LB2D_shift_2 ) : ( n120 ) ;
assign n122 =  ( n37 ) ? ( LB2D_shift_3 ) : ( LB2D_shift_3 ) ;
assign n123 =  ( n32 ) ? ( LB2D_shift_3 ) : ( n122 ) ;
assign n124 =  ( n25 ) ? ( LB2D_shift_2 ) : ( n123 ) ;
assign n125 =  ( n18 ) ? ( LB2D_shift_3 ) : ( n124 ) ;
assign n126 =  ( n9 ) ? ( LB2D_shift_3 ) : ( n125 ) ;
assign n127 =  ( n4 ) ? ( LB2D_shift_3 ) : ( n126 ) ;
assign n128 =  ( n37 ) ? ( LB2D_shift_4 ) : ( LB2D_shift_4 ) ;
assign n129 =  ( n32 ) ? ( LB2D_shift_4 ) : ( n128 ) ;
assign n130 =  ( n25 ) ? ( LB2D_shift_3 ) : ( n129 ) ;
assign n131 =  ( n18 ) ? ( LB2D_shift_4 ) : ( n130 ) ;
assign n132 =  ( n9 ) ? ( LB2D_shift_4 ) : ( n131 ) ;
assign n133 =  ( n4 ) ? ( LB2D_shift_4 ) : ( n132 ) ;
assign n134 =  ( n37 ) ? ( LB2D_shift_5 ) : ( LB2D_shift_5 ) ;
assign n135 =  ( n32 ) ? ( LB2D_shift_5 ) : ( n134 ) ;
assign n136 =  ( n25 ) ? ( LB2D_shift_4 ) : ( n135 ) ;
assign n137 =  ( n18 ) ? ( LB2D_shift_5 ) : ( n136 ) ;
assign n138 =  ( n9 ) ? ( LB2D_shift_5 ) : ( n137 ) ;
assign n139 =  ( n4 ) ? ( LB2D_shift_5 ) : ( n138 ) ;
assign n140 =  ( n37 ) ? ( LB2D_shift_6 ) : ( LB2D_shift_6 ) ;
assign n141 =  ( n32 ) ? ( LB2D_shift_6 ) : ( n140 ) ;
assign n142 =  ( n25 ) ? ( LB2D_shift_5 ) : ( n141 ) ;
assign n143 =  ( n18 ) ? ( LB2D_shift_6 ) : ( n142 ) ;
assign n144 =  ( n9 ) ? ( LB2D_shift_6 ) : ( n143 ) ;
assign n145 =  ( n4 ) ? ( LB2D_shift_6 ) : ( n144 ) ;
assign n146 =  ( n37 ) ? ( LB2D_shift_7 ) : ( LB2D_shift_7 ) ;
assign n147 =  ( n32 ) ? ( LB2D_shift_7 ) : ( n146 ) ;
assign n148 =  ( n25 ) ? ( LB2D_shift_6 ) : ( n147 ) ;
assign n149 =  ( n18 ) ? ( LB2D_shift_7 ) : ( n148 ) ;
assign n150 =  ( n9 ) ? ( LB2D_shift_7 ) : ( n149 ) ;
assign n151 =  ( n4 ) ? ( LB2D_shift_7 ) : ( n150 ) ;
assign n152 =  ( LB2D_shift_x ) + ( 9'd1 )  ;
assign n153 =  ( n37 ) ? ( LB2D_shift_x ) : ( LB2D_shift_x ) ;
assign n154 =  ( n32 ) ? ( LB2D_shift_x ) : ( n153 ) ;
assign n155 =  ( n25 ) ? ( n152 ) : ( n154 ) ;
assign n156 =  ( n18 ) ? ( LB2D_shift_x ) : ( n155 ) ;
assign n157 =  ( n9 ) ? ( LB2D_shift_x ) : ( n156 ) ;
assign n158 =  ( n4 ) ? ( LB2D_shift_x ) : ( n157 ) ;
assign n159 =  ( LB2D_shift_y ) < ( 10'd480 )  ;
assign n160 =  ( LB2D_shift_x ) < ( 9'd488 )  ;
assign n161 =  ( LB2D_shift_y ) + ( 10'd1 )  ;
assign n162 =  ( n160 ) ? ( LB2D_shift_y ) : ( n161 ) ;
assign n163 =  ( n159 ) ? ( n162 ) : ( 10'd480 ) ;
assign n164 =  ( n37 ) ? ( LB2D_shift_y ) : ( LB2D_shift_y ) ;
assign n165 =  ( n32 ) ? ( LB2D_shift_y ) : ( n164 ) ;
assign n166 =  ( n25 ) ? ( n163 ) : ( n165 ) ;
assign n167 =  ( n18 ) ? ( LB2D_shift_y ) : ( n166 ) ;
assign n168 =  ( n9 ) ? ( LB2D_shift_y ) : ( n167 ) ;
assign n169 =  ( n4 ) ? ( LB2D_shift_y ) : ( n168 ) ;
assign n170 =  ( stencil_stream_full ) == ( 1'd1 )  ;
assign n171 =  ( n170 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_0 ) ;
assign n172 = gb_fun(n171) ;
assign n173 =  ( n37 ) ? ( arg_0_TDATA ) : ( arg_0_TDATA ) ;
assign n174 =  ( n32 ) ? ( arg_0_TDATA ) : ( n173 ) ;
assign n175 =  ( n25 ) ? ( arg_0_TDATA ) : ( n174 ) ;
assign n176 =  ( n18 ) ? ( n172 ) : ( n175 ) ;
assign n177 =  ( n9 ) ? ( arg_0_TDATA ) : ( n176 ) ;
assign n178 =  ( n4 ) ? ( arg_0_TDATA ) : ( n177 ) ;
assign n179 =  ( gb_pp_it_8 ) == ( 1'd1 )  ;
assign n180 =  ( n179 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n181 =  ( n37 ) ? ( arg_0_TVALID ) : ( arg_0_TVALID ) ;
assign n182 =  ( n32 ) ? ( arg_0_TVALID ) : ( n181 ) ;
assign n183 =  ( n25 ) ? ( arg_0_TVALID ) : ( n182 ) ;
assign n184 =  ( n18 ) ? ( n180 ) : ( n183 ) ;
assign n185 =  ( n9 ) ? ( arg_0_TVALID ) : ( n184 ) ;
assign n186 =  ( n4 ) ? ( 1'd0 ) : ( n185 ) ;
assign n187 =  ( n37 ) ? ( 1'd1 ) : ( arg_1_TREADY ) ;
assign n188 =  ( n51 ) ? ( 1'd1 ) : ( n187 ) ;
assign n189 =  ( n32 ) ? ( arg_1_TREADY ) : ( n188 ) ;
assign n190 =  ( n25 ) ? ( arg_1_TREADY ) : ( n189 ) ;
assign n191 =  ( n18 ) ? ( arg_1_TREADY ) : ( n190 ) ;
assign n192 =  ( n9 ) ? ( 1'd0 ) : ( n191 ) ;
assign n193 =  ( n4 ) ? ( 1'd0 ) : ( n192 ) ;
assign n194 =  ( gb_p_cnt ) + ( 19'd1 )  ;
assign n195 =  ( n194 ) == ( 19'd307200 )  ;
assign n196 =  ( n195 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n197 =  ( n37 ) ? ( gb_exit_it_1 ) : ( gb_exit_it_1 ) ;
assign n198 =  ( n32 ) ? ( gb_exit_it_1 ) : ( n197 ) ;
assign n199 =  ( n25 ) ? ( gb_exit_it_1 ) : ( n198 ) ;
assign n200 =  ( n18 ) ? ( n196 ) : ( n199 ) ;
assign n201 =  ( n9 ) ? ( gb_exit_it_1 ) : ( n200 ) ;
assign n202 =  ( n4 ) ? ( gb_exit_it_1 ) : ( n201 ) ;
assign n203 =  ( n37 ) ? ( gb_exit_it_2 ) : ( gb_exit_it_2 ) ;
assign n204 =  ( n32 ) ? ( gb_exit_it_2 ) : ( n203 ) ;
assign n205 =  ( n25 ) ? ( gb_exit_it_2 ) : ( n204 ) ;
assign n206 =  ( n18 ) ? ( gb_exit_it_1 ) : ( n205 ) ;
assign n207 =  ( n9 ) ? ( gb_exit_it_2 ) : ( n206 ) ;
assign n208 =  ( n4 ) ? ( gb_exit_it_2 ) : ( n207 ) ;
assign n209 =  ( n37 ) ? ( gb_exit_it_3 ) : ( gb_exit_it_3 ) ;
assign n210 =  ( n32 ) ? ( gb_exit_it_3 ) : ( n209 ) ;
assign n211 =  ( n25 ) ? ( gb_exit_it_3 ) : ( n210 ) ;
assign n212 =  ( n18 ) ? ( gb_exit_it_2 ) : ( n211 ) ;
assign n213 =  ( n9 ) ? ( gb_exit_it_3 ) : ( n212 ) ;
assign n214 =  ( n4 ) ? ( gb_exit_it_3 ) : ( n213 ) ;
assign n215 =  ( n37 ) ? ( gb_exit_it_4 ) : ( gb_exit_it_4 ) ;
assign n216 =  ( n32 ) ? ( gb_exit_it_4 ) : ( n215 ) ;
assign n217 =  ( n25 ) ? ( gb_exit_it_4 ) : ( n216 ) ;
assign n218 =  ( n18 ) ? ( gb_exit_it_3 ) : ( n217 ) ;
assign n219 =  ( n9 ) ? ( gb_exit_it_4 ) : ( n218 ) ;
assign n220 =  ( n4 ) ? ( gb_exit_it_4 ) : ( n219 ) ;
assign n221 =  ( n37 ) ? ( gb_exit_it_5 ) : ( gb_exit_it_5 ) ;
assign n222 =  ( n32 ) ? ( gb_exit_it_5 ) : ( n221 ) ;
assign n223 =  ( n25 ) ? ( gb_exit_it_5 ) : ( n222 ) ;
assign n224 =  ( n18 ) ? ( gb_exit_it_4 ) : ( n223 ) ;
assign n225 =  ( n9 ) ? ( gb_exit_it_5 ) : ( n224 ) ;
assign n226 =  ( n4 ) ? ( gb_exit_it_5 ) : ( n225 ) ;
assign n227 =  ( n37 ) ? ( gb_exit_it_6 ) : ( gb_exit_it_6 ) ;
assign n228 =  ( n32 ) ? ( gb_exit_it_6 ) : ( n227 ) ;
assign n229 =  ( n25 ) ? ( gb_exit_it_6 ) : ( n228 ) ;
assign n230 =  ( n18 ) ? ( gb_exit_it_5 ) : ( n229 ) ;
assign n231 =  ( n9 ) ? ( gb_exit_it_6 ) : ( n230 ) ;
assign n232 =  ( n4 ) ? ( gb_exit_it_6 ) : ( n231 ) ;
assign n233 =  ( n37 ) ? ( gb_exit_it_7 ) : ( gb_exit_it_7 ) ;
assign n234 =  ( n32 ) ? ( gb_exit_it_7 ) : ( n233 ) ;
assign n235 =  ( n25 ) ? ( gb_exit_it_7 ) : ( n234 ) ;
assign n236 =  ( n18 ) ? ( gb_exit_it_6 ) : ( n235 ) ;
assign n237 =  ( n9 ) ? ( gb_exit_it_7 ) : ( n236 ) ;
assign n238 =  ( n4 ) ? ( gb_exit_it_7 ) : ( n237 ) ;
assign n239 =  ( n37 ) ? ( gb_exit_it_8 ) : ( gb_exit_it_8 ) ;
assign n240 =  ( n32 ) ? ( gb_exit_it_8 ) : ( n239 ) ;
assign n241 =  ( n25 ) ? ( gb_exit_it_8 ) : ( n240 ) ;
assign n242 =  ( n18 ) ? ( gb_exit_it_7 ) : ( n241 ) ;
assign n243 =  ( n9 ) ? ( gb_exit_it_8 ) : ( n242 ) ;
assign n244 =  ( n4 ) ? ( gb_exit_it_8 ) : ( n243 ) ;
assign n245 =  ( gb_p_cnt ) < ( 19'd307200 )  ;
assign n246 =  ( n245 ) ? ( n194 ) : ( 19'd307200 ) ;
assign n247 =  ( n37 ) ? ( gb_p_cnt ) : ( gb_p_cnt ) ;
assign n248 =  ( n32 ) ? ( gb_p_cnt ) : ( n247 ) ;
assign n249 =  ( n25 ) ? ( gb_p_cnt ) : ( n248 ) ;
assign n250 =  ( n18 ) ? ( n246 ) : ( n249 ) ;
assign n251 =  ( n9 ) ? ( gb_p_cnt ) : ( n250 ) ;
assign n252 =  ( n4 ) ? ( gb_p_cnt ) : ( n251 ) ;
assign n253 =  ( n37 ) ? ( gb_pp_it_1 ) : ( gb_pp_it_1 ) ;
assign n254 =  ( n32 ) ? ( gb_pp_it_1 ) : ( n253 ) ;
assign n255 =  ( n25 ) ? ( gb_pp_it_1 ) : ( n254 ) ;
assign n256 =  ( n18 ) ? ( 1'd1 ) : ( n255 ) ;
assign n257 =  ( n9 ) ? ( gb_pp_it_1 ) : ( n256 ) ;
assign n258 =  ( n4 ) ? ( gb_pp_it_1 ) : ( n257 ) ;
assign n259 =  ( n37 ) ? ( gb_pp_it_2 ) : ( gb_pp_it_2 ) ;
assign n260 =  ( n32 ) ? ( gb_pp_it_2 ) : ( n259 ) ;
assign n261 =  ( n25 ) ? ( gb_pp_it_2 ) : ( n260 ) ;
assign n262 =  ( n18 ) ? ( gb_pp_it_1 ) : ( n261 ) ;
assign n263 =  ( n9 ) ? ( gb_pp_it_2 ) : ( n262 ) ;
assign n264 =  ( n4 ) ? ( gb_pp_it_2 ) : ( n263 ) ;
assign n265 =  ( n37 ) ? ( gb_pp_it_3 ) : ( gb_pp_it_3 ) ;
assign n266 =  ( n32 ) ? ( gb_pp_it_3 ) : ( n265 ) ;
assign n267 =  ( n25 ) ? ( gb_pp_it_3 ) : ( n266 ) ;
assign n268 =  ( n18 ) ? ( gb_pp_it_2 ) : ( n267 ) ;
assign n269 =  ( n9 ) ? ( gb_pp_it_3 ) : ( n268 ) ;
assign n270 =  ( n4 ) ? ( gb_pp_it_3 ) : ( n269 ) ;
assign n271 =  ( n37 ) ? ( gb_pp_it_4 ) : ( gb_pp_it_4 ) ;
assign n272 =  ( n32 ) ? ( gb_pp_it_4 ) : ( n271 ) ;
assign n273 =  ( n25 ) ? ( gb_pp_it_4 ) : ( n272 ) ;
assign n274 =  ( n18 ) ? ( gb_pp_it_3 ) : ( n273 ) ;
assign n275 =  ( n9 ) ? ( gb_pp_it_4 ) : ( n274 ) ;
assign n276 =  ( n4 ) ? ( gb_pp_it_4 ) : ( n275 ) ;
assign n277 =  ( n37 ) ? ( gb_pp_it_5 ) : ( gb_pp_it_5 ) ;
assign n278 =  ( n32 ) ? ( gb_pp_it_5 ) : ( n277 ) ;
assign n279 =  ( n25 ) ? ( gb_pp_it_5 ) : ( n278 ) ;
assign n280 =  ( n18 ) ? ( gb_pp_it_4 ) : ( n279 ) ;
assign n281 =  ( n9 ) ? ( gb_pp_it_5 ) : ( n280 ) ;
assign n282 =  ( n4 ) ? ( gb_pp_it_5 ) : ( n281 ) ;
assign n283 =  ( n37 ) ? ( gb_pp_it_6 ) : ( gb_pp_it_6 ) ;
assign n284 =  ( n32 ) ? ( gb_pp_it_6 ) : ( n283 ) ;
assign n285 =  ( n25 ) ? ( gb_pp_it_6 ) : ( n284 ) ;
assign n286 =  ( n18 ) ? ( gb_pp_it_5 ) : ( n285 ) ;
assign n287 =  ( n9 ) ? ( gb_pp_it_6 ) : ( n286 ) ;
assign n288 =  ( n4 ) ? ( gb_pp_it_6 ) : ( n287 ) ;
assign n289 =  ( n37 ) ? ( gb_pp_it_7 ) : ( gb_pp_it_7 ) ;
assign n290 =  ( n32 ) ? ( gb_pp_it_7 ) : ( n289 ) ;
assign n291 =  ( n25 ) ? ( gb_pp_it_7 ) : ( n290 ) ;
assign n292 =  ( n18 ) ? ( gb_pp_it_6 ) : ( n291 ) ;
assign n293 =  ( n9 ) ? ( gb_pp_it_7 ) : ( n292 ) ;
assign n294 =  ( n4 ) ? ( gb_pp_it_7 ) : ( n293 ) ;
assign n295 =  ( n37 ) ? ( gb_pp_it_8 ) : ( gb_pp_it_8 ) ;
assign n296 =  ( n32 ) ? ( gb_pp_it_8 ) : ( n295 ) ;
assign n297 =  ( n25 ) ? ( gb_pp_it_8 ) : ( n296 ) ;
assign n298 =  ( n18 ) ? ( gb_pp_it_7 ) : ( n297 ) ;
assign n299 =  ( n9 ) ? ( gb_pp_it_8 ) : ( n298 ) ;
assign n300 =  ( n4 ) ? ( gb_pp_it_8 ) : ( n299 ) ;
assign n301 =  ( n37 ) ? ( gb_pp_it_9 ) : ( gb_pp_it_9 ) ;
assign n302 =  ( n32 ) ? ( gb_pp_it_9 ) : ( n301 ) ;
assign n303 =  ( n25 ) ? ( gb_pp_it_9 ) : ( n302 ) ;
assign n304 =  ( n18 ) ? ( gb_pp_it_8 ) : ( n303 ) ;
assign n305 =  ( n9 ) ? ( gb_pp_it_9 ) : ( n304 ) ;
assign n306 =  ( n4 ) ? ( gb_pp_it_9 ) : ( n305 ) ;
assign n307 =  ( n37 ) ? ( LB1D_buff ) : ( in_stream_buff_0 ) ;
assign n308 =  ( n32 ) ? ( in_stream_buff_0 ) : ( n307 ) ;
assign n309 =  ( n25 ) ? ( in_stream_buff_0 ) : ( n308 ) ;
assign n310 =  ( n18 ) ? ( in_stream_buff_0 ) : ( n309 ) ;
assign n311 =  ( n9 ) ? ( in_stream_buff_0 ) : ( n310 ) ;
assign n312 =  ( n4 ) ? ( in_stream_buff_0 ) : ( n311 ) ;
assign n313 =  ( n37 ) ? ( in_stream_buff_0 ) : ( in_stream_buff_1 ) ;
assign n314 =  ( n32 ) ? ( in_stream_buff_1 ) : ( n313 ) ;
assign n315 =  ( n25 ) ? ( in_stream_buff_1 ) : ( n314 ) ;
assign n316 =  ( n18 ) ? ( in_stream_buff_1 ) : ( n315 ) ;
assign n317 =  ( n9 ) ? ( in_stream_buff_1 ) : ( n316 ) ;
assign n318 =  ( n4 ) ? ( in_stream_buff_1 ) : ( n317 ) ;
assign n319 =  ( in_stream_full ) == ( 1'd1 )  ;
assign n320 =  ( n319 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n321 =  ( n37 ) ? ( 1'd0 ) : ( in_stream_empty ) ;
assign n322 =  ( n32 ) ? ( n320 ) : ( n321 ) ;
assign n323 =  ( n25 ) ? ( in_stream_empty ) : ( n322 ) ;
assign n324 =  ( n18 ) ? ( in_stream_empty ) : ( n323 ) ;
assign n325 =  ( n9 ) ? ( in_stream_empty ) : ( n324 ) ;
assign n326 =  ( n4 ) ? ( in_stream_empty ) : ( n325 ) ;
assign n327 =  ( in_stream_empty ) == ( 1'd1 )  ;
assign n328 =  ( n327 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n329 =  ( n37 ) ? ( n328 ) : ( in_stream_full ) ;
assign n330 =  ( n32 ) ? ( 1'd0 ) : ( n329 ) ;
assign n331 =  ( n25 ) ? ( in_stream_full ) : ( n330 ) ;
assign n332 =  ( n18 ) ? ( in_stream_full ) : ( n331 ) ;
assign n333 =  ( n9 ) ? ( in_stream_full ) : ( n332 ) ;
assign n334 =  ( n4 ) ? ( in_stream_full ) : ( n333 ) ;
assign n335 =  ( n319 ) ? ( in_stream_buff_1 ) : ( in_stream_buff_0 ) ;
assign n336 =  ( LB2D_proc_w ) == ( 64'd0 )  ;
assign n337 =  (  LB2D_proc_7 [ LB2D_proc_x ] )  ;
assign n338 =  ( LB2D_proc_w ) == ( 64'd1 )  ;
assign n339 =  (  LB2D_proc_0 [ LB2D_proc_x ] )  ;
assign n340 =  ( LB2D_proc_w ) == ( 64'd2 )  ;
assign n341 =  (  LB2D_proc_1 [ LB2D_proc_x ] )  ;
assign n342 =  ( LB2D_proc_w ) == ( 64'd3 )  ;
assign n343 =  (  LB2D_proc_2 [ LB2D_proc_x ] )  ;
assign n344 =  ( LB2D_proc_w ) == ( 64'd4 )  ;
assign n345 =  (  LB2D_proc_3 [ LB2D_proc_x ] )  ;
assign n346 =  ( LB2D_proc_w ) == ( 64'd5 )  ;
assign n347 =  (  LB2D_proc_4 [ LB2D_proc_x ] )  ;
assign n348 =  ( LB2D_proc_w ) == ( 64'd6 )  ;
assign n349 =  (  LB2D_proc_5 [ LB2D_proc_x ] )  ;
assign n350 =  (  LB2D_proc_6 [ LB2D_proc_x ] )  ;
assign n351 =  ( n348 ) ? ( n349 ) : ( n350 ) ;
assign n352 =  ( n346 ) ? ( n347 ) : ( n351 ) ;
assign n353 =  ( n344 ) ? ( n345 ) : ( n352 ) ;
assign n354 =  ( n342 ) ? ( n343 ) : ( n353 ) ;
assign n355 =  ( n340 ) ? ( n341 ) : ( n354 ) ;
assign n356 =  ( n338 ) ? ( n339 ) : ( n355 ) ;
assign n357 =  ( n336 ) ? ( n337 ) : ( n356 ) ;
assign n358 =  ( n348 ) ? ( n347 ) : ( n349 ) ;
assign n359 =  ( n346 ) ? ( n345 ) : ( n358 ) ;
assign n360 =  ( n344 ) ? ( n343 ) : ( n359 ) ;
assign n361 =  ( n342 ) ? ( n341 ) : ( n360 ) ;
assign n362 =  ( n340 ) ? ( n339 ) : ( n361 ) ;
assign n363 =  ( n338 ) ? ( n337 ) : ( n362 ) ;
assign n364 =  ( n336 ) ? ( n350 ) : ( n363 ) ;
assign n365 =  ( n348 ) ? ( n345 ) : ( n347 ) ;
assign n366 =  ( n346 ) ? ( n343 ) : ( n365 ) ;
assign n367 =  ( n344 ) ? ( n341 ) : ( n366 ) ;
assign n368 =  ( n342 ) ? ( n339 ) : ( n367 ) ;
assign n369 =  ( n340 ) ? ( n337 ) : ( n368 ) ;
assign n370 =  ( n338 ) ? ( n350 ) : ( n369 ) ;
assign n371 =  ( n336 ) ? ( n349 ) : ( n370 ) ;
assign n372 =  ( n348 ) ? ( n343 ) : ( n345 ) ;
assign n373 =  ( n346 ) ? ( n341 ) : ( n372 ) ;
assign n374 =  ( n344 ) ? ( n339 ) : ( n373 ) ;
assign n375 =  ( n342 ) ? ( n337 ) : ( n374 ) ;
assign n376 =  ( n340 ) ? ( n350 ) : ( n375 ) ;
assign n377 =  ( n338 ) ? ( n349 ) : ( n376 ) ;
assign n378 =  ( n336 ) ? ( n347 ) : ( n377 ) ;
assign n379 =  ( n348 ) ? ( n341 ) : ( n343 ) ;
assign n380 =  ( n346 ) ? ( n339 ) : ( n379 ) ;
assign n381 =  ( n344 ) ? ( n337 ) : ( n380 ) ;
assign n382 =  ( n342 ) ? ( n350 ) : ( n381 ) ;
assign n383 =  ( n340 ) ? ( n349 ) : ( n382 ) ;
assign n384 =  ( n338 ) ? ( n347 ) : ( n383 ) ;
assign n385 =  ( n336 ) ? ( n345 ) : ( n384 ) ;
assign n386 =  ( n348 ) ? ( n339 ) : ( n341 ) ;
assign n387 =  ( n346 ) ? ( n337 ) : ( n386 ) ;
assign n388 =  ( n344 ) ? ( n350 ) : ( n387 ) ;
assign n389 =  ( n342 ) ? ( n349 ) : ( n388 ) ;
assign n390 =  ( n340 ) ? ( n347 ) : ( n389 ) ;
assign n391 =  ( n338 ) ? ( n345 ) : ( n390 ) ;
assign n392 =  ( n336 ) ? ( n343 ) : ( n391 ) ;
assign n393 =  ( n348 ) ? ( n337 ) : ( n339 ) ;
assign n394 =  ( n346 ) ? ( n350 ) : ( n393 ) ;
assign n395 =  ( n344 ) ? ( n349 ) : ( n394 ) ;
assign n396 =  ( n342 ) ? ( n347 ) : ( n395 ) ;
assign n397 =  ( n340 ) ? ( n345 ) : ( n396 ) ;
assign n398 =  ( n338 ) ? ( n343 ) : ( n397 ) ;
assign n399 =  ( n336 ) ? ( n341 ) : ( n398 ) ;
assign n400 =  ( n348 ) ? ( n350 ) : ( n337 ) ;
assign n401 =  ( n346 ) ? ( n349 ) : ( n400 ) ;
assign n402 =  ( n344 ) ? ( n347 ) : ( n401 ) ;
assign n403 =  ( n342 ) ? ( n345 ) : ( n402 ) ;
assign n404 =  ( n340 ) ? ( n343 ) : ( n403 ) ;
assign n405 =  ( n338 ) ? ( n341 ) : ( n404 ) ;
assign n406 =  ( n336 ) ? ( n339 ) : ( n405 ) ;
assign n407 =  { ( n399 ) , ( n406 ) }  ;
assign n408 =  { ( n392 ) , ( n407 ) }  ;
assign n409 =  { ( n385 ) , ( n408 ) }  ;
assign n410 =  { ( n378 ) , ( n409 ) }  ;
assign n411 =  { ( n371 ) , ( n410 ) }  ;
assign n412 =  { ( n364 ) , ( n411 ) }  ;
assign n413 =  { ( n357 ) , ( n412 ) }  ;
assign n414 =  { ( n335 ) , ( n413 ) }  ;
assign n415 =  ( n30 ) ? ( slice_stream_buff_0 ) : ( n414 ) ;
assign n416 =  ( n37 ) ? ( slice_stream_buff_0 ) : ( slice_stream_buff_0 ) ;
assign n417 =  ( n32 ) ? ( n415 ) : ( n416 ) ;
assign n418 =  ( n25 ) ? ( slice_stream_buff_0 ) : ( n417 ) ;
assign n419 =  ( n18 ) ? ( slice_stream_buff_0 ) : ( n418 ) ;
assign n420 =  ( n9 ) ? ( slice_stream_buff_0 ) : ( n419 ) ;
assign n421 =  ( n4 ) ? ( slice_stream_buff_0 ) : ( n420 ) ;
assign n422 =  ( n30 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n423 =  ( n37 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_1 ) ;
assign n424 =  ( n32 ) ? ( n422 ) : ( n423 ) ;
assign n425 =  ( n25 ) ? ( slice_stream_buff_1 ) : ( n424 ) ;
assign n426 =  ( n18 ) ? ( slice_stream_buff_1 ) : ( n425 ) ;
assign n427 =  ( n9 ) ? ( slice_stream_buff_1 ) : ( n426 ) ;
assign n428 =  ( n4 ) ? ( slice_stream_buff_1 ) : ( n427 ) ;
assign n429 =  ( n102 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n430 =  ( n30 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n431 =  ( n37 ) ? ( slice_stream_empty ) : ( slice_stream_empty ) ;
assign n432 =  ( n32 ) ? ( n430 ) : ( n431 ) ;
assign n433 =  ( n25 ) ? ( n429 ) : ( n432 ) ;
assign n434 =  ( n18 ) ? ( slice_stream_empty ) : ( n433 ) ;
assign n435 =  ( n9 ) ? ( slice_stream_empty ) : ( n434 ) ;
assign n436 =  ( n4 ) ? ( slice_stream_empty ) : ( n435 ) ;
assign n437 =  ( slice_stream_empty ) == ( 1'd1 )  ;
assign n438 =  ( n437 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n439 =  ( n30 ) ? ( 1'd0 ) : ( n438 ) ;
assign n440 =  ( n37 ) ? ( slice_stream_full ) : ( slice_stream_full ) ;
assign n441 =  ( n32 ) ? ( n439 ) : ( n440 ) ;
assign n442 =  ( n25 ) ? ( 1'd0 ) : ( n441 ) ;
assign n443 =  ( n18 ) ? ( slice_stream_full ) : ( n442 ) ;
assign n444 =  ( n9 ) ? ( slice_stream_full ) : ( n443 ) ;
assign n445 =  ( n4 ) ? ( slice_stream_full ) : ( n444 ) ;
assign n446 =  ( LB2D_shift_x ) >= ( 9'd8 )  ;
assign n447 = n103[71:64] ;
assign n448 = LB2D_shift_0[71:64] ;
assign n449 = LB2D_shift_1[71:64] ;
assign n450 = LB2D_shift_2[71:64] ;
assign n451 = LB2D_shift_3[71:64] ;
assign n452 = LB2D_shift_4[71:64] ;
assign n453 = LB2D_shift_5[71:64] ;
assign n454 = LB2D_shift_6[71:64] ;
assign n455 = LB2D_shift_7[71:64] ;
assign n456 =  { ( n454 ) , ( n455 ) }  ;
assign n457 =  { ( n453 ) , ( n456 ) }  ;
assign n458 =  { ( n452 ) , ( n457 ) }  ;
assign n459 =  { ( n451 ) , ( n458 ) }  ;
assign n460 =  { ( n450 ) , ( n459 ) }  ;
assign n461 =  { ( n449 ) , ( n460 ) }  ;
assign n462 =  { ( n448 ) , ( n461 ) }  ;
assign n463 =  { ( n447 ) , ( n462 ) }  ;
assign n464 = n103[63:56] ;
assign n465 = LB2D_shift_0[63:56] ;
assign n466 = LB2D_shift_1[63:56] ;
assign n467 = LB2D_shift_2[63:56] ;
assign n468 = LB2D_shift_3[63:56] ;
assign n469 = LB2D_shift_4[63:56] ;
assign n470 = LB2D_shift_5[63:56] ;
assign n471 = LB2D_shift_6[63:56] ;
assign n472 = LB2D_shift_7[63:56] ;
assign n473 =  { ( n471 ) , ( n472 ) }  ;
assign n474 =  { ( n470 ) , ( n473 ) }  ;
assign n475 =  { ( n469 ) , ( n474 ) }  ;
assign n476 =  { ( n468 ) , ( n475 ) }  ;
assign n477 =  { ( n467 ) , ( n476 ) }  ;
assign n478 =  { ( n466 ) , ( n477 ) }  ;
assign n479 =  { ( n465 ) , ( n478 ) }  ;
assign n480 =  { ( n464 ) , ( n479 ) }  ;
assign n481 = n103[55:48] ;
assign n482 = LB2D_shift_0[55:48] ;
assign n483 = LB2D_shift_1[55:48] ;
assign n484 = LB2D_shift_2[55:48] ;
assign n485 = LB2D_shift_3[55:48] ;
assign n486 = LB2D_shift_4[55:48] ;
assign n487 = LB2D_shift_5[55:48] ;
assign n488 = LB2D_shift_6[55:48] ;
assign n489 = LB2D_shift_7[55:48] ;
assign n490 =  { ( n488 ) , ( n489 ) }  ;
assign n491 =  { ( n487 ) , ( n490 ) }  ;
assign n492 =  { ( n486 ) , ( n491 ) }  ;
assign n493 =  { ( n485 ) , ( n492 ) }  ;
assign n494 =  { ( n484 ) , ( n493 ) }  ;
assign n495 =  { ( n483 ) , ( n494 ) }  ;
assign n496 =  { ( n482 ) , ( n495 ) }  ;
assign n497 =  { ( n481 ) , ( n496 ) }  ;
assign n498 = n103[47:40] ;
assign n499 = LB2D_shift_0[47:40] ;
assign n500 = LB2D_shift_1[47:40] ;
assign n501 = LB2D_shift_2[47:40] ;
assign n502 = LB2D_shift_3[47:40] ;
assign n503 = LB2D_shift_4[47:40] ;
assign n504 = LB2D_shift_5[47:40] ;
assign n505 = LB2D_shift_6[47:40] ;
assign n506 = LB2D_shift_7[47:40] ;
assign n507 =  { ( n505 ) , ( n506 ) }  ;
assign n508 =  { ( n504 ) , ( n507 ) }  ;
assign n509 =  { ( n503 ) , ( n508 ) }  ;
assign n510 =  { ( n502 ) , ( n509 ) }  ;
assign n511 =  { ( n501 ) , ( n510 ) }  ;
assign n512 =  { ( n500 ) , ( n511 ) }  ;
assign n513 =  { ( n499 ) , ( n512 ) }  ;
assign n514 =  { ( n498 ) , ( n513 ) }  ;
assign n515 = n103[39:32] ;
assign n516 = LB2D_shift_0[39:32] ;
assign n517 = LB2D_shift_1[39:32] ;
assign n518 = LB2D_shift_2[39:32] ;
assign n519 = LB2D_shift_3[39:32] ;
assign n520 = LB2D_shift_4[39:32] ;
assign n521 = LB2D_shift_5[39:32] ;
assign n522 = LB2D_shift_6[39:32] ;
assign n523 = LB2D_shift_7[39:32] ;
assign n524 =  { ( n522 ) , ( n523 ) }  ;
assign n525 =  { ( n521 ) , ( n524 ) }  ;
assign n526 =  { ( n520 ) , ( n525 ) }  ;
assign n527 =  { ( n519 ) , ( n526 ) }  ;
assign n528 =  { ( n518 ) , ( n527 ) }  ;
assign n529 =  { ( n517 ) , ( n528 ) }  ;
assign n530 =  { ( n516 ) , ( n529 ) }  ;
assign n531 =  { ( n515 ) , ( n530 ) }  ;
assign n532 = n103[31:24] ;
assign n533 = LB2D_shift_0[31:24] ;
assign n534 = LB2D_shift_1[31:24] ;
assign n535 = LB2D_shift_2[31:24] ;
assign n536 = LB2D_shift_3[31:24] ;
assign n537 = LB2D_shift_4[31:24] ;
assign n538 = LB2D_shift_5[31:24] ;
assign n539 = LB2D_shift_6[31:24] ;
assign n540 = LB2D_shift_7[31:24] ;
assign n541 =  { ( n539 ) , ( n540 ) }  ;
assign n542 =  { ( n538 ) , ( n541 ) }  ;
assign n543 =  { ( n537 ) , ( n542 ) }  ;
assign n544 =  { ( n536 ) , ( n543 ) }  ;
assign n545 =  { ( n535 ) , ( n544 ) }  ;
assign n546 =  { ( n534 ) , ( n545 ) }  ;
assign n547 =  { ( n533 ) , ( n546 ) }  ;
assign n548 =  { ( n532 ) , ( n547 ) }  ;
assign n549 = n103[23:16] ;
assign n550 = LB2D_shift_0[23:16] ;
assign n551 = LB2D_shift_1[23:16] ;
assign n552 = LB2D_shift_2[23:16] ;
assign n553 = LB2D_shift_3[23:16] ;
assign n554 = LB2D_shift_4[23:16] ;
assign n555 = LB2D_shift_5[23:16] ;
assign n556 = LB2D_shift_6[23:16] ;
assign n557 = LB2D_shift_7[23:16] ;
assign n558 =  { ( n556 ) , ( n557 ) }  ;
assign n559 =  { ( n555 ) , ( n558 ) }  ;
assign n560 =  { ( n554 ) , ( n559 ) }  ;
assign n561 =  { ( n553 ) , ( n560 ) }  ;
assign n562 =  { ( n552 ) , ( n561 ) }  ;
assign n563 =  { ( n551 ) , ( n562 ) }  ;
assign n564 =  { ( n550 ) , ( n563 ) }  ;
assign n565 =  { ( n549 ) , ( n564 ) }  ;
assign n566 = n103[15:8] ;
assign n567 = LB2D_shift_0[15:8] ;
assign n568 = LB2D_shift_1[15:8] ;
assign n569 = LB2D_shift_2[15:8] ;
assign n570 = LB2D_shift_3[15:8] ;
assign n571 = LB2D_shift_4[15:8] ;
assign n572 = LB2D_shift_5[15:8] ;
assign n573 = LB2D_shift_6[15:8] ;
assign n574 = LB2D_shift_7[15:8] ;
assign n575 =  { ( n573 ) , ( n574 ) }  ;
assign n576 =  { ( n572 ) , ( n575 ) }  ;
assign n577 =  { ( n571 ) , ( n576 ) }  ;
assign n578 =  { ( n570 ) , ( n577 ) }  ;
assign n579 =  { ( n569 ) , ( n578 ) }  ;
assign n580 =  { ( n568 ) , ( n579 ) }  ;
assign n581 =  { ( n567 ) , ( n580 ) }  ;
assign n582 =  { ( n566 ) , ( n581 ) }  ;
assign n583 = n103[7:0] ;
assign n584 = LB2D_shift_0[7:0] ;
assign n585 = LB2D_shift_1[7:0] ;
assign n586 = LB2D_shift_2[7:0] ;
assign n587 = LB2D_shift_3[7:0] ;
assign n588 = LB2D_shift_4[7:0] ;
assign n589 = LB2D_shift_5[7:0] ;
assign n590 = LB2D_shift_6[7:0] ;
assign n591 = LB2D_shift_7[7:0] ;
assign n592 =  { ( n590 ) , ( n591 ) }  ;
assign n593 =  { ( n589 ) , ( n592 ) }  ;
assign n594 =  { ( n588 ) , ( n593 ) }  ;
assign n595 =  { ( n587 ) , ( n594 ) }  ;
assign n596 =  { ( n586 ) , ( n595 ) }  ;
assign n597 =  { ( n585 ) , ( n596 ) }  ;
assign n598 =  { ( n584 ) , ( n597 ) }  ;
assign n599 =  { ( n583 ) , ( n598 ) }  ;
assign n600 =  { ( n582 ) , ( n599 ) }  ;
assign n601 =  { ( n565 ) , ( n600 ) }  ;
assign n602 =  { ( n548 ) , ( n601 ) }  ;
assign n603 =  { ( n531 ) , ( n602 ) }  ;
assign n604 =  { ( n514 ) , ( n603 ) }  ;
assign n605 =  { ( n497 ) , ( n604 ) }  ;
assign n606 =  { ( n480 ) , ( n605 ) }  ;
assign n607 =  { ( n463 ) , ( n606 ) }  ;
assign n608 =  ( n446 ) ? ( n607 ) : ( stencil_stream_buff_0 ) ;
assign n609 =  ( n37 ) ? ( stencil_stream_buff_0 ) : ( stencil_stream_buff_0 ) ;
assign n610 =  ( n32 ) ? ( stencil_stream_buff_0 ) : ( n609 ) ;
assign n611 =  ( n25 ) ? ( n608 ) : ( n610 ) ;
assign n612 =  ( n18 ) ? ( stencil_stream_buff_0 ) : ( n611 ) ;
assign n613 =  ( n9 ) ? ( stencil_stream_buff_0 ) : ( n612 ) ;
assign n614 =  ( n4 ) ? ( stencil_stream_buff_0 ) : ( n613 ) ;
assign n615 =  ( n37 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_1 ) ;
assign n616 =  ( n32 ) ? ( stencil_stream_buff_1 ) : ( n615 ) ;
assign n617 =  ( n25 ) ? ( stencil_stream_buff_0 ) : ( n616 ) ;
assign n618 =  ( n18 ) ? ( stencil_stream_buff_1 ) : ( n617 ) ;
assign n619 =  ( n9 ) ? ( stencil_stream_buff_1 ) : ( n618 ) ;
assign n620 =  ( n4 ) ? ( stencil_stream_buff_1 ) : ( n619 ) ;
assign n621 =  ( n170 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n622 =  ( n23 ) ? ( stencil_stream_empty ) : ( 1'd0 ) ;
assign n623 =  ( n37 ) ? ( stencil_stream_empty ) : ( stencil_stream_empty ) ;
assign n624 =  ( n32 ) ? ( stencil_stream_empty ) : ( n623 ) ;
assign n625 =  ( n25 ) ? ( n622 ) : ( n624 ) ;
assign n626 =  ( n18 ) ? ( n621 ) : ( n625 ) ;
assign n627 =  ( n9 ) ? ( stencil_stream_empty ) : ( n626 ) ;
assign n628 =  ( n4 ) ? ( stencil_stream_empty ) : ( n627 ) ;
assign n629 =  ( n14 ) ? ( 1'd0 ) : ( 1'd0 ) ;
assign n630 =  ( stencil_stream_empty ) == ( 1'd1 )  ;
assign n631 =  ( n630 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n632 =  ( n23 ) ? ( stencil_stream_full ) : ( n631 ) ;
assign n633 =  ( n37 ) ? ( stencil_stream_full ) : ( stencil_stream_full ) ;
assign n634 =  ( n32 ) ? ( stencil_stream_full ) : ( n633 ) ;
assign n635 =  ( n25 ) ? ( n632 ) : ( n634 ) ;
assign n636 =  ( n18 ) ? ( n629 ) : ( n635 ) ;
assign n637 =  ( n9 ) ? ( stencil_stream_full ) : ( n636 ) ;
assign n638 =  ( n4 ) ? ( stencil_stream_full ) : ( n637 ) ;
assign n639 = ~ ( n4 ) ;
assign n640 = ~ ( n9 ) ;
assign n641 =  ( n639 ) & ( n640 )  ;
assign n642 = ~ ( n18 ) ;
assign n643 =  ( n641 ) & ( n642 )  ;
assign n644 = ~ ( n25 ) ;
assign n645 =  ( n643 ) & ( n644 )  ;
assign n646 = ~ ( n32 ) ;
assign n647 =  ( n645 ) & ( n646 )  ;
assign n648 = ~ ( n37 ) ;
assign n649 =  ( n647 ) & ( n648 )  ;
assign n650 =  ( n647 ) & ( n37 )  ;
assign n651 =  ( n645 ) & ( n32 )  ;
assign n652 = ~ ( n336 ) ;
assign n653 =  ( n651 ) & ( n652 )  ;
assign n654 =  ( n651 ) & ( n336 )  ;
assign n655 =  ( n643 ) & ( n25 )  ;
assign n656 =  ( n641 ) & ( n18 )  ;
assign n657 =  ( n639 ) & ( n9 )  ;
assign LB2D_proc_0_addr0 = n654 ? (LB2D_proc_x) : (0);
assign LB2D_proc_0_data0 = n654 ? (n335) : (LB2D_proc_0[0]);
assign n658 = ~ ( n338 ) ;
assign n659 =  ( n651 ) & ( n658 )  ;
assign n660 =  ( n651 ) & ( n338 )  ;
assign LB2D_proc_1_addr0 = n660 ? (LB2D_proc_x) : (0);
assign LB2D_proc_1_data0 = n660 ? (n335) : (LB2D_proc_1[0]);
assign n661 = ~ ( n340 ) ;
assign n662 =  ( n651 ) & ( n661 )  ;
assign n663 =  ( n651 ) & ( n340 )  ;
assign LB2D_proc_2_addr0 = n663 ? (LB2D_proc_x) : (0);
assign LB2D_proc_2_data0 = n663 ? (n335) : (LB2D_proc_2[0]);
assign n664 = ~ ( n342 ) ;
assign n665 =  ( n651 ) & ( n664 )  ;
assign n666 =  ( n651 ) & ( n342 )  ;
assign LB2D_proc_3_addr0 = n666 ? (LB2D_proc_x) : (0);
assign LB2D_proc_3_data0 = n666 ? (n335) : (LB2D_proc_3[0]);
assign n667 = ~ ( n344 ) ;
assign n668 =  ( n651 ) & ( n667 )  ;
assign n669 =  ( n651 ) & ( n344 )  ;
assign LB2D_proc_4_addr0 = n669 ? (LB2D_proc_x) : (0);
assign LB2D_proc_4_data0 = n669 ? (n335) : (LB2D_proc_4[0]);
assign n670 = ~ ( n346 ) ;
assign n671 =  ( n651 ) & ( n670 )  ;
assign n672 =  ( n651 ) & ( n346 )  ;
assign LB2D_proc_5_addr0 = n672 ? (LB2D_proc_x) : (0);
assign LB2D_proc_5_data0 = n672 ? (n335) : (LB2D_proc_5[0]);
assign n673 = ~ ( n348 ) ;
assign n674 =  ( n651 ) & ( n673 )  ;
assign n675 =  ( n651 ) & ( n348 )  ;
assign LB2D_proc_6_addr0 = n675 ? (LB2D_proc_x) : (0);
assign LB2D_proc_6_data0 = n675 ? (n335) : (LB2D_proc_6[0]);
assign n676 = ~ ( n72 ) ;
assign n677 =  ( n651 ) & ( n676 )  ;
assign n678 =  ( n651 ) & ( n72 )  ;
assign LB2D_proc_7_addr0 = n678 ? (LB2D_proc_x) : (0);
assign LB2D_proc_7_data0 = n678 ? (n335) : (LB2D_proc_7[0]);
function [7:0] gb_fun ;
input [647:0] arg0;
    begin
//TODO: Add the specific function HERE.    end
endfunction

always @(posedge clk) begin
   if(rst) begin
       LB1D_buff <= LB1D_buff;
       LB1D_in <= LB1D_in;
       LB1D_it_1 <= LB1D_it_1;
       LB1D_p_cnt <= LB1D_p_cnt;
       LB1D_uIn <= LB1D_uIn;
       LB2D_proc_w <= LB2D_proc_w;
       LB2D_proc_x <= LB2D_proc_x;
       LB2D_proc_y <= LB2D_proc_y;
       LB2D_shift_0 <= LB2D_shift_0;
       LB2D_shift_1 <= LB2D_shift_1;
       LB2D_shift_2 <= LB2D_shift_2;
       LB2D_shift_3 <= LB2D_shift_3;
       LB2D_shift_4 <= LB2D_shift_4;
       LB2D_shift_5 <= LB2D_shift_5;
       LB2D_shift_6 <= LB2D_shift_6;
       LB2D_shift_7 <= LB2D_shift_7;
       LB2D_shift_x <= LB2D_shift_x;
       LB2D_shift_y <= LB2D_shift_y;
       arg_0_TDATA <= arg_0_TDATA;
       arg_0_TVALID <= arg_0_TVALID;
       arg_1_TREADY <= arg_1_TREADY;
       gb_exit_it_1 <= gb_exit_it_1;
       gb_exit_it_2 <= gb_exit_it_2;
       gb_exit_it_3 <= gb_exit_it_3;
       gb_exit_it_4 <= gb_exit_it_4;
       gb_exit_it_5 <= gb_exit_it_5;
       gb_exit_it_6 <= gb_exit_it_6;
       gb_exit_it_7 <= gb_exit_it_7;
       gb_exit_it_8 <= gb_exit_it_8;
       gb_p_cnt <= gb_p_cnt;
       gb_pp_it_1 <= gb_pp_it_1;
       gb_pp_it_2 <= gb_pp_it_2;
       gb_pp_it_3 <= gb_pp_it_3;
       gb_pp_it_4 <= gb_pp_it_4;
       gb_pp_it_5 <= gb_pp_it_5;
       gb_pp_it_6 <= gb_pp_it_6;
       gb_pp_it_7 <= gb_pp_it_7;
       gb_pp_it_8 <= gb_pp_it_8;
       gb_pp_it_9 <= gb_pp_it_9;
       in_stream_buff_0 <= in_stream_buff_0;
       in_stream_buff_1 <= in_stream_buff_1;
       in_stream_empty <= in_stream_empty;
       in_stream_full <= in_stream_full;
       slice_stream_buff_0 <= slice_stream_buff_0;
       slice_stream_buff_1 <= slice_stream_buff_1;
       slice_stream_empty <= slice_stream_empty;
       slice_stream_full <= slice_stream_full;
       stencil_stream_buff_0 <= stencil_stream_buff_0;
       stencil_stream_buff_1 <= stencil_stream_buff_1;
       stencil_stream_empty <= stencil_stream_empty;
       stencil_stream_full <= stencil_stream_full;
   end
   else if(step) begin
       LB1D_buff <= n43;
       LB1D_in <= n49;
       LB1D_it_1 <= n52;
       LB1D_p_cnt <= n63;
       LB1D_uIn <= n68;
       LB2D_proc_w <= n81;
       LB2D_proc_x <= n91;
       LB2D_proc_y <= n101;
       LB2D_shift_0 <= n109;
       LB2D_shift_1 <= n115;
       LB2D_shift_2 <= n121;
       LB2D_shift_3 <= n127;
       LB2D_shift_4 <= n133;
       LB2D_shift_5 <= n139;
       LB2D_shift_6 <= n145;
       LB2D_shift_7 <= n151;
       LB2D_shift_x <= n158;
       LB2D_shift_y <= n169;
       arg_0_TDATA <= n178;
       arg_0_TVALID <= n186;
       arg_1_TREADY <= n193;
       gb_exit_it_1 <= n202;
       gb_exit_it_2 <= n208;
       gb_exit_it_3 <= n214;
       gb_exit_it_4 <= n220;
       gb_exit_it_5 <= n226;
       gb_exit_it_6 <= n232;
       gb_exit_it_7 <= n238;
       gb_exit_it_8 <= n244;
       gb_p_cnt <= n252;
       gb_pp_it_1 <= n258;
       gb_pp_it_2 <= n264;
       gb_pp_it_3 <= n270;
       gb_pp_it_4 <= n276;
       gb_pp_it_5 <= n282;
       gb_pp_it_6 <= n288;
       gb_pp_it_7 <= n294;
       gb_pp_it_8 <= n300;
       gb_pp_it_9 <= n306;
       in_stream_buff_0 <= n312;
       in_stream_buff_1 <= n318;
       in_stream_empty <= n326;
       in_stream_full <= n334;
       slice_stream_buff_0 <= n421;
       slice_stream_buff_1 <= n428;
       slice_stream_empty <= n436;
       slice_stream_full <= n445;
       stencil_stream_buff_0 <= n614;
       stencil_stream_buff_1 <= n620;
       stencil_stream_empty <= n628;
       stencil_stream_full <= n638;
       LB2D_proc_0 [ LB2D_proc_0_addr0 ] <= LB2D_proc_0_data0;
       LB2D_proc_1 [ LB2D_proc_1_addr0 ] <= LB2D_proc_1_data0;
       LB2D_proc_2 [ LB2D_proc_2_addr0 ] <= LB2D_proc_2_data0;
       LB2D_proc_3 [ LB2D_proc_3_addr0 ] <= LB2D_proc_3_data0;
       LB2D_proc_4 [ LB2D_proc_4_addr0 ] <= LB2D_proc_4_data0;
       LB2D_proc_5 [ LB2D_proc_5_addr0 ] <= LB2D_proc_5_data0;
       LB2D_proc_6 [ LB2D_proc_6_addr0 ] <= LB2D_proc_6_data0;
       LB2D_proc_7 [ LB2D_proc_7_addr0 ] <= LB2D_proc_7_data0;
   end
end
endmodule
