module GB(
arg_0_TREADY,
arg_1_TDATA,
arg_1_TVALID,
LB1D_buff,
LB2D_proc_w,
LB2D_proc_x,
LB2D_proc_y,
LB2D_shift_0,
LB2D_shift_1,
LB2D_shift_2,
LB2D_shift_3,
LB2D_shift_4,
LB2D_shift_5,
LB2D_shift_6,
LB2D_shift_7,
LB2D_shift_x,
LB2D_shift_y,
arg_0_TDATA,
arg_0_TVALID,
arg_1_TREADY,
gb_exit_it_1,
gb_exit_it_2,
gb_exit_it_3,
gb_exit_it_4,
gb_exit_it_5,
gb_exit_it_6,
gb_exit_it_7,
gb_exit_it_8,
gb_pp_it_1,
gb_pp_it_2,
gb_pp_it_3,
gb_pp_it_4,
gb_pp_it_5,
gb_pp_it_6,
gb_pp_it_7,
gb_pp_it_8,
gb_pp_it_9,
in_stream_buff_0,
in_stream_buff_1,
in_stream_empty,
in_stream_full,
p_cnt,
slice_stream_buff_0,
slice_stream_buff_1,
slice_stream_empty,
slice_stream_full,
stencil_stream_buff_0,
stencil_stream_buff_1,
stencil_stream_empty,
stencil_stream_full,
clk,rst,
step
);
input            arg_0_TREADY;
input      [7:0] arg_1_TDATA;
input            arg_1_TVALID;
input clk;
input rst;
input step;
output      [7:0] LB1D_buff;
output     [63:0] LB2D_proc_w;
output      [8:0] LB2D_proc_x;
output      [9:0] LB2D_proc_y;
output     [71:0] LB2D_shift_0;
output     [71:0] LB2D_shift_1;
output     [71:0] LB2D_shift_2;
output     [71:0] LB2D_shift_3;
output     [71:0] LB2D_shift_4;
output     [71:0] LB2D_shift_5;
output     [71:0] LB2D_shift_6;
output     [71:0] LB2D_shift_7;
output      [8:0] LB2D_shift_x;
output      [9:0] LB2D_shift_y;
output      [7:0] arg_0_TDATA;
output            arg_0_TVALID;
output            arg_1_TREADY;
output            gb_exit_it_1;
output            gb_exit_it_2;
output            gb_exit_it_3;
output            gb_exit_it_4;
output            gb_exit_it_5;
output            gb_exit_it_6;
output            gb_exit_it_7;
output            gb_exit_it_8;
output            gb_pp_it_1;
output            gb_pp_it_2;
output            gb_pp_it_3;
output            gb_pp_it_4;
output            gb_pp_it_5;
output            gb_pp_it_6;
output            gb_pp_it_7;
output            gb_pp_it_8;
output            gb_pp_it_9;
output      [7:0] in_stream_buff_0;
output      [7:0] in_stream_buff_1;
output            in_stream_empty;
output            in_stream_full;
output     [18:0] p_cnt;
output     [71:0] slice_stream_buff_0;
output     [71:0] slice_stream_buff_1;
output            slice_stream_empty;
output            slice_stream_full;
output    [647:0] stencil_stream_buff_0;
output    [647:0] stencil_stream_buff_1;
output            stencil_stream_empty;
output            stencil_stream_full;
reg      [7:0] LB1D_buff;
reg     [63:0] LB2D_proc_w;
reg      [8:0] LB2D_proc_x;
reg      [9:0] LB2D_proc_y;
reg     [71:0] LB2D_shift_0;
reg     [71:0] LB2D_shift_1;
reg     [71:0] LB2D_shift_2;
reg     [71:0] LB2D_shift_3;
reg     [71:0] LB2D_shift_4;
reg     [71:0] LB2D_shift_5;
reg     [71:0] LB2D_shift_6;
reg     [71:0] LB2D_shift_7;
reg      [8:0] LB2D_shift_x;
reg      [9:0] LB2D_shift_y;
reg      [7:0] arg_0_TDATA;
reg            arg_0_TVALID;
reg            arg_1_TREADY;
reg            gb_exit_it_1;
reg            gb_exit_it_2;
reg            gb_exit_it_3;
reg            gb_exit_it_4;
reg            gb_exit_it_5;
reg            gb_exit_it_6;
reg            gb_exit_it_7;
reg            gb_exit_it_8;
reg            gb_pp_it_1;
reg            gb_pp_it_2;
reg            gb_pp_it_3;
reg            gb_pp_it_4;
reg            gb_pp_it_5;
reg            gb_pp_it_6;
reg            gb_pp_it_7;
reg            gb_pp_it_8;
reg            gb_pp_it_9;
reg      [7:0] in_stream_buff_0;
reg      [7:0] in_stream_buff_1;
reg            in_stream_empty;
reg            in_stream_full;
reg     [18:0] p_cnt;
reg     [71:0] slice_stream_buff_0;
reg     [71:0] slice_stream_buff_1;
reg            slice_stream_empty;
reg            slice_stream_full;
reg    [647:0] stencil_stream_buff_0;
reg    [647:0] stencil_stream_buff_1;
reg            stencil_stream_empty;
reg            stencil_stream_full;
wire            arg_0_TREADY;
wire      [7:0] arg_1_TDATA;
wire            arg_1_TVALID;
wire            n0;
wire            n1;
wire            n2;
wire            n3;
wire            n4;
wire            n5;
wire            n6;
wire            n7;
wire            n8;
wire            n9;
wire            n10;
wire            n11;
wire            n12;
wire            n13;
wire            n14;
wire            n15;
wire            n16;
wire            n17;
wire            n18;
wire            n19;
wire            n20;
wire            n21;
wire            n22;
wire            n23;
wire            n24;
wire            n25;
wire            n26;
wire            n27;
wire            n28;
wire            n29;
wire            n30;
wire            n31;
wire      [7:0] n32;
wire      [7:0] n33;
wire      [7:0] n34;
wire      [7:0] n35;
wire      [7:0] n36;
wire      [7:0] n37;
wire            n38;
wire            n39;
wire     [63:0] n40;
wire     [63:0] n41;
wire     [63:0] n42;
wire     [63:0] n43;
wire     [63:0] n44;
wire     [63:0] n45;
wire     [63:0] n46;
wire     [63:0] n47;
wire     [63:0] n48;
wire      [8:0] n49;
wire      [8:0] n50;
wire      [8:0] n51;
wire      [8:0] n52;
wire      [8:0] n53;
wire      [8:0] n54;
wire      [8:0] n55;
wire      [8:0] n56;
wire            n57;
wire      [9:0] n58;
wire      [9:0] n59;
wire      [9:0] n60;
wire      [9:0] n61;
wire      [9:0] n62;
wire      [9:0] n63;
wire      [9:0] n64;
wire      [9:0] n65;
wire      [9:0] n66;
wire            n67;
wire     [71:0] n68;
wire     [71:0] n69;
wire     [71:0] n70;
wire     [71:0] n71;
wire     [71:0] n72;
wire     [71:0] n73;
wire     [71:0] n74;
wire     [71:0] n75;
wire     [71:0] n76;
wire     [71:0] n77;
wire     [71:0] n78;
wire     [71:0] n79;
wire     [71:0] n80;
wire     [71:0] n81;
wire     [71:0] n82;
wire     [71:0] n83;
wire     [71:0] n84;
wire     [71:0] n85;
wire     [71:0] n86;
wire     [71:0] n87;
wire     [71:0] n88;
wire     [71:0] n89;
wire     [71:0] n90;
wire     [71:0] n91;
wire     [71:0] n92;
wire     [71:0] n93;
wire     [71:0] n94;
wire     [71:0] n95;
wire     [71:0] n96;
wire     [71:0] n97;
wire     [71:0] n98;
wire     [71:0] n99;
wire     [71:0] n100;
wire     [71:0] n101;
wire     [71:0] n102;
wire     [71:0] n103;
wire     [71:0] n104;
wire     [71:0] n105;
wire     [71:0] n106;
wire     [71:0] n107;
wire     [71:0] n108;
wire     [71:0] n109;
wire     [71:0] n110;
wire     [71:0] n111;
wire     [71:0] n112;
wire     [71:0] n113;
wire     [71:0] n114;
wire     [71:0] n115;
wire     [71:0] n116;
wire            n117;
wire      [8:0] n118;
wire      [8:0] n119;
wire      [8:0] n120;
wire      [8:0] n121;
wire      [8:0] n122;
wire      [8:0] n123;
wire      [8:0] n124;
wire      [8:0] n125;
wire            n126;
wire      [9:0] n127;
wire      [9:0] n128;
wire      [9:0] n129;
wire      [9:0] n130;
wire      [9:0] n131;
wire      [9:0] n132;
wire      [9:0] n133;
wire      [9:0] n134;
wire      [9:0] n135;
wire            n136;
wire    [647:0] n137;
wire      [7:0] n138;
wire      [7:0] n139;
wire      [7:0] n140;
wire      [7:0] n141;
wire      [7:0] n142;
wire      [7:0] n143;
wire      [7:0] n144;
wire            n145;
wire            n146;
wire            n147;
wire            n148;
wire            n149;
wire            n150;
wire            n151;
wire            n152;
wire            n153;
wire            n154;
wire            n155;
wire            n156;
wire            n157;
wire            n158;
wire     [18:0] n159;
wire            n160;
wire            n161;
wire            n162;
wire            n163;
wire            n164;
wire            n165;
wire            n166;
wire            n167;
wire            n168;
wire            n169;
wire            n170;
wire            n171;
wire            n172;
wire            n173;
wire            n174;
wire            n175;
wire            n176;
wire            n177;
wire            n178;
wire      [7:0] n179;
wire      [7:0] n180;
wire      [7:0] n181;
wire      [7:0] n182;
wire      [7:0] n183;
wire      [7:0] n184;
wire      [7:0] n185;
wire      [7:0] n186;
wire      [7:0] n187;
wire      [7:0] n188;
wire      [7:0] n189;
wire      [7:0] n190;
wire            n191;
wire            n192;
wire            n193;
wire            n194;
wire            n195;
wire            n196;
wire            n197;
wire            n198;
wire            n199;
wire            n200;
wire            n201;
wire            n202;
wire            n203;
wire            n204;
wire            n205;
wire            n206;
wire            n207;
wire     [18:0] n208;
wire     [18:0] n209;
wire      [7:0] n210;
wire            n211;
wire      [7:0] n212;
wire            n213;
wire      [7:0] n214;
wire            n215;
wire      [7:0] n216;
wire            n217;
wire      [7:0] n218;
wire            n219;
wire      [7:0] n220;
wire            n221;
wire      [7:0] n222;
wire            n223;
wire      [7:0] n224;
wire      [7:0] n225;
wire      [7:0] n226;
wire      [7:0] n227;
wire      [7:0] n228;
wire      [7:0] n229;
wire      [7:0] n230;
wire      [7:0] n231;
wire      [7:0] n232;
wire      [7:0] n233;
wire      [7:0] n234;
wire      [7:0] n235;
wire      [7:0] n236;
wire      [7:0] n237;
wire      [7:0] n238;
wire      [7:0] n239;
wire      [7:0] n240;
wire      [7:0] n241;
wire      [7:0] n242;
wire      [7:0] n243;
wire      [7:0] n244;
wire      [7:0] n245;
wire      [7:0] n246;
wire      [7:0] n247;
wire      [7:0] n248;
wire      [7:0] n249;
wire      [7:0] n250;
wire      [7:0] n251;
wire      [7:0] n252;
wire      [7:0] n253;
wire      [7:0] n254;
wire      [7:0] n255;
wire      [7:0] n256;
wire      [7:0] n257;
wire      [7:0] n258;
wire      [7:0] n259;
wire      [7:0] n260;
wire      [7:0] n261;
wire      [7:0] n262;
wire      [7:0] n263;
wire      [7:0] n264;
wire      [7:0] n265;
wire      [7:0] n266;
wire      [7:0] n267;
wire      [7:0] n268;
wire      [7:0] n269;
wire      [7:0] n270;
wire      [7:0] n271;
wire      [7:0] n272;
wire      [7:0] n273;
wire      [7:0] n274;
wire      [7:0] n275;
wire      [7:0] n276;
wire      [7:0] n277;
wire      [7:0] n278;
wire      [7:0] n279;
wire      [7:0] n280;
wire      [7:0] n281;
wire     [15:0] n282;
wire     [23:0] n283;
wire     [31:0] n284;
wire     [39:0] n285;
wire     [47:0] n286;
wire     [55:0] n287;
wire     [63:0] n288;
wire     [71:0] n289;
wire     [71:0] n290;
wire     [71:0] n291;
wire     [71:0] n292;
wire     [71:0] n293;
wire     [71:0] n294;
wire     [71:0] n295;
wire     [71:0] n296;
wire     [71:0] n297;
wire     [71:0] n298;
wire     [71:0] n299;
wire     [71:0] n300;
wire     [71:0] n301;
wire     [71:0] n302;
wire     [71:0] n303;
wire            n304;
wire            n305;
wire            n306;
wire            n307;
wire            n308;
wire            n309;
wire            n310;
wire            n311;
wire            n312;
wire            n313;
wire            n314;
wire            n315;
wire            n316;
wire            n317;
wire            n318;
wire            n319;
wire            n320;
wire            n321;
wire      [7:0] n322;
wire      [7:0] n323;
wire      [7:0] n324;
wire      [7:0] n325;
wire      [7:0] n326;
wire      [7:0] n327;
wire      [7:0] n328;
wire      [7:0] n329;
wire      [7:0] n330;
wire     [15:0] n331;
wire     [23:0] n332;
wire     [31:0] n333;
wire     [39:0] n334;
wire     [47:0] n335;
wire     [55:0] n336;
wire     [63:0] n337;
wire     [71:0] n338;
wire      [7:0] n339;
wire      [7:0] n340;
wire      [7:0] n341;
wire      [7:0] n342;
wire      [7:0] n343;
wire      [7:0] n344;
wire      [7:0] n345;
wire      [7:0] n346;
wire      [7:0] n347;
wire     [15:0] n348;
wire     [23:0] n349;
wire     [31:0] n350;
wire     [39:0] n351;
wire     [47:0] n352;
wire     [55:0] n353;
wire     [63:0] n354;
wire     [71:0] n355;
wire      [7:0] n356;
wire      [7:0] n357;
wire      [7:0] n358;
wire      [7:0] n359;
wire      [7:0] n360;
wire      [7:0] n361;
wire      [7:0] n362;
wire      [7:0] n363;
wire      [7:0] n364;
wire     [15:0] n365;
wire     [23:0] n366;
wire     [31:0] n367;
wire     [39:0] n368;
wire     [47:0] n369;
wire     [55:0] n370;
wire     [63:0] n371;
wire     [71:0] n372;
wire      [7:0] n373;
wire      [7:0] n374;
wire      [7:0] n375;
wire      [7:0] n376;
wire      [7:0] n377;
wire      [7:0] n378;
wire      [7:0] n379;
wire      [7:0] n380;
wire      [7:0] n381;
wire     [15:0] n382;
wire     [23:0] n383;
wire     [31:0] n384;
wire     [39:0] n385;
wire     [47:0] n386;
wire     [55:0] n387;
wire     [63:0] n388;
wire     [71:0] n389;
wire      [7:0] n390;
wire      [7:0] n391;
wire      [7:0] n392;
wire      [7:0] n393;
wire      [7:0] n394;
wire      [7:0] n395;
wire      [7:0] n396;
wire      [7:0] n397;
wire      [7:0] n398;
wire     [15:0] n399;
wire     [23:0] n400;
wire     [31:0] n401;
wire     [39:0] n402;
wire     [47:0] n403;
wire     [55:0] n404;
wire     [63:0] n405;
wire     [71:0] n406;
wire      [7:0] n407;
wire      [7:0] n408;
wire      [7:0] n409;
wire      [7:0] n410;
wire      [7:0] n411;
wire      [7:0] n412;
wire      [7:0] n413;
wire      [7:0] n414;
wire      [7:0] n415;
wire     [15:0] n416;
wire     [23:0] n417;
wire     [31:0] n418;
wire     [39:0] n419;
wire     [47:0] n420;
wire     [55:0] n421;
wire     [63:0] n422;
wire     [71:0] n423;
wire      [7:0] n424;
wire      [7:0] n425;
wire      [7:0] n426;
wire      [7:0] n427;
wire      [7:0] n428;
wire      [7:0] n429;
wire      [7:0] n430;
wire      [7:0] n431;
wire      [7:0] n432;
wire     [15:0] n433;
wire     [23:0] n434;
wire     [31:0] n435;
wire     [39:0] n436;
wire     [47:0] n437;
wire     [55:0] n438;
wire     [63:0] n439;
wire     [71:0] n440;
wire      [7:0] n441;
wire      [7:0] n442;
wire      [7:0] n443;
wire      [7:0] n444;
wire      [7:0] n445;
wire      [7:0] n446;
wire      [7:0] n447;
wire      [7:0] n448;
wire      [7:0] n449;
wire     [15:0] n450;
wire     [23:0] n451;
wire     [31:0] n452;
wire     [39:0] n453;
wire     [47:0] n454;
wire     [55:0] n455;
wire     [63:0] n456;
wire     [71:0] n457;
wire      [7:0] n458;
wire      [7:0] n459;
wire      [7:0] n460;
wire      [7:0] n461;
wire      [7:0] n462;
wire      [7:0] n463;
wire      [7:0] n464;
wire      [7:0] n465;
wire      [7:0] n466;
wire     [15:0] n467;
wire     [23:0] n468;
wire     [31:0] n469;
wire     [39:0] n470;
wire     [47:0] n471;
wire     [55:0] n472;
wire     [63:0] n473;
wire     [71:0] n474;
wire    [143:0] n475;
wire    [215:0] n476;
wire    [287:0] n477;
wire    [359:0] n478;
wire    [431:0] n479;
wire    [503:0] n480;
wire    [575:0] n481;
wire    [647:0] n482;
wire    [647:0] n483;
wire    [647:0] n484;
wire    [647:0] n485;
wire    [647:0] n486;
wire    [647:0] n487;
wire    [647:0] n488;
wire    [647:0] n489;
wire    [647:0] n490;
wire    [647:0] n491;
wire    [647:0] n492;
wire    [647:0] n493;
wire    [647:0] n494;
wire    [647:0] n495;
wire            n496;
wire            n497;
wire            n498;
wire            n499;
wire            n500;
wire            n501;
wire            n502;
wire            n503;
wire            n504;
wire            n505;
wire            n506;
wire            n507;
wire            n508;
wire            n509;
wire            n510;
wire            n511;
wire            n512;
wire            n513;
wire      [8:0] LB2D_proc_0_addr0;
wire      [7:0] LB2D_proc_0_data0;
wire            n514;
wire            n515;
wire            n516;
wire            n517;
wire            n518;
wire            n519;
wire            n520;
wire            n521;
wire            n522;
wire            n523;
wire            n524;
wire            n525;
wire            n526;
wire            n527;
wire            n528;
wire            n529;
wire            n530;
wire            n531;
wire            n532;
wire      [8:0] LB2D_proc_1_addr0;
wire      [7:0] LB2D_proc_1_data0;
wire            n533;
wire            n534;
wire            n535;
wire      [8:0] LB2D_proc_2_addr0;
wire      [7:0] LB2D_proc_2_data0;
wire            n536;
wire            n537;
wire            n538;
wire      [8:0] LB2D_proc_3_addr0;
wire      [7:0] LB2D_proc_3_data0;
wire            n539;
wire            n540;
wire            n541;
wire      [8:0] LB2D_proc_4_addr0;
wire      [7:0] LB2D_proc_4_data0;
wire            n542;
wire            n543;
wire            n544;
wire      [8:0] LB2D_proc_5_addr0;
wire      [7:0] LB2D_proc_5_data0;
wire            n545;
wire            n546;
wire            n547;
wire      [8:0] LB2D_proc_6_addr0;
wire      [7:0] LB2D_proc_6_data0;
wire            n548;
wire            n549;
wire            n550;
wire      [8:0] LB2D_proc_7_addr0;
wire      [7:0] LB2D_proc_7_data0;
wire            n551;
wire            n552;
wire            n553;
wire            n554;
reg      [7:0] LB2D_proc_0[511:0];
reg      [7:0] LB2D_proc_1[511:0];
reg      [7:0] LB2D_proc_2[511:0];
reg      [7:0] LB2D_proc_3[511:0];
reg      [7:0] LB2D_proc_4[511:0];
reg      [7:0] LB2D_proc_5[511:0];
reg      [7:0] LB2D_proc_6[511:0];
reg      [7:0] LB2D_proc_7[511:0];
wire clk;
wire rst;
wire step;
assign n0 =  ( arg_0_TREADY ) == ( 1'd1 )  ;
assign n1 =  ( arg_0_TVALID ) == ( 1'd1 )  ;
assign n2 =  ( n0 ) & ( n1 )  ;
assign n3 =  ( arg_1_TVALID ) == ( 1'd0 )  ;
assign n4 =  ( n2 ) & ( n3 )  ;
assign n5 =  ( arg_1_TREADY ) == ( 1'd1 )  ;
assign n6 =  ( arg_1_TVALID ) == ( 1'd1 )  ;
assign n7 =  ( n5 ) & ( n6 )  ;
assign n8 =  ( arg_0_TREADY ) == ( 1'd0 )  ;
assign n9 =  ( n7 ) & ( n8 )  ;
assign n10 =  ( arg_0_TVALID ) == ( 1'd0 )  ;
assign n11 =  ( gb_exit_it_1 ) == ( 1'd0 )  ;
assign n12 =  ( stencil_stream_empty ) == ( 1'd0 )  ;
assign n13 =  ( n11 ) & ( n12 )  ;
assign n14 =  ( gb_exit_it_1 ) == ( 1'd1 )  ;
assign n15 =  ( gb_exit_it_8 ) == ( 1'd0 )  ;
assign n16 =  ( n14 ) & ( n15 )  ;
assign n17 =  ( n13 ) | ( n16 )  ;
assign n18 =  ( n10 ) & ( n17 )  ;
assign n19 =  ( slice_stream_empty ) == ( 1'd0 )  ;
assign n20 =  ( stencil_stream_full ) == ( 1'd0 )  ;
assign n21 =  ( LB2D_shift_x ) < ( 9'd8 )  ;
assign n22 =  ( n20 ) | ( n21 )  ;
assign n23 =  ( n19 ) & ( n22 )  ;
assign n24 =  ( in_stream_empty ) == ( 1'd0 )  ;
assign n25 =  ( slice_stream_full ) == ( 1'd0 )  ;
assign n26 =  ( LB2D_proc_y ) < ( 10'd8 )  ;
assign n27 =  ( n25 ) | ( n26 )  ;
assign n28 =  ( n24 ) & ( n27 )  ;
assign n29 =  ( arg_1_TREADY ) == ( 1'd0 )  ;
assign n30 =  ( in_stream_full ) == ( 1'd0 )  ;
assign n31 =  ( n29 ) & ( n30 )  ;
assign n32 =  ( n31 ) ? ( LB1D_buff ) : ( LB1D_buff ) ;
assign n33 =  ( n28 ) ? ( LB1D_buff ) : ( n32 ) ;
assign n34 =  ( n23 ) ? ( LB1D_buff ) : ( n33 ) ;
assign n35 =  ( n18 ) ? ( LB1D_buff ) : ( n34 ) ;
assign n36 =  ( n9 ) ? ( arg_1_TDATA ) : ( n35 ) ;
assign n37 =  ( n4 ) ? ( arg_1_TDATA ) : ( n36 ) ;
assign n38 =  ( LB2D_proc_w ) < ( 64'd7 )  ;
assign n39 =  ( LB2D_proc_x ) < ( 9'd487 )  ;
assign n40 =  ( LB2D_proc_w ) + ( 64'd1 )  ;
assign n41 =  ( n39 ) ? ( LB2D_proc_w ) : ( n40 ) ;
assign n42 =  ( n38 ) ? ( n41 ) : ( 64'd0 ) ;
assign n43 =  ( n31 ) ? ( LB2D_proc_w ) : ( LB2D_proc_w ) ;
assign n44 =  ( n28 ) ? ( n42 ) : ( n43 ) ;
assign n45 =  ( n23 ) ? ( LB2D_proc_w ) : ( n44 ) ;
assign n46 =  ( n18 ) ? ( LB2D_proc_w ) : ( n45 ) ;
assign n47 =  ( n9 ) ? ( LB2D_proc_w ) : ( n46 ) ;
assign n48 =  ( n4 ) ? ( LB2D_proc_w ) : ( n47 ) ;
assign n49 =  ( LB2D_proc_x ) + ( 9'd1 )  ;
assign n50 =  ( n39 ) ? ( n49 ) : ( 9'd0 ) ;
assign n51 =  ( n31 ) ? ( LB2D_proc_x ) : ( LB2D_proc_x ) ;
assign n52 =  ( n28 ) ? ( n50 ) : ( n51 ) ;
assign n53 =  ( n23 ) ? ( LB2D_proc_x ) : ( n52 ) ;
assign n54 =  ( n18 ) ? ( LB2D_proc_x ) : ( n53 ) ;
assign n55 =  ( n9 ) ? ( LB2D_proc_x ) : ( n54 ) ;
assign n56 =  ( n4 ) ? ( LB2D_proc_x ) : ( n55 ) ;
assign n57 =  ( LB2D_proc_y ) < ( 10'd487 )  ;
assign n58 =  ( LB2D_proc_y ) + ( 10'd1 )  ;
assign n59 =  ( n39 ) ? ( LB2D_proc_y ) : ( n58 ) ;
assign n60 =  ( n57 ) ? ( n59 ) : ( 10'd487 ) ;
assign n61 =  ( n31 ) ? ( LB2D_proc_y ) : ( LB2D_proc_y ) ;
assign n62 =  ( n28 ) ? ( n60 ) : ( n61 ) ;
assign n63 =  ( n23 ) ? ( LB2D_proc_y ) : ( n62 ) ;
assign n64 =  ( n18 ) ? ( LB2D_proc_y ) : ( n63 ) ;
assign n65 =  ( n9 ) ? ( LB2D_proc_y ) : ( n64 ) ;
assign n66 =  ( n4 ) ? ( LB2D_proc_y ) : ( n65 ) ;
assign n67 =  ( slice_stream_full ) == ( 1'd1 )  ;
assign n68 =  ( n67 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n69 =  ( n31 ) ? ( LB2D_shift_0 ) : ( LB2D_shift_0 ) ;
assign n70 =  ( n28 ) ? ( LB2D_shift_0 ) : ( n69 ) ;
assign n71 =  ( n23 ) ? ( n68 ) : ( n70 ) ;
assign n72 =  ( n18 ) ? ( LB2D_shift_0 ) : ( n71 ) ;
assign n73 =  ( n9 ) ? ( LB2D_shift_0 ) : ( n72 ) ;
assign n74 =  ( n4 ) ? ( LB2D_shift_0 ) : ( n73 ) ;
assign n75 =  ( n31 ) ? ( LB2D_shift_1 ) : ( LB2D_shift_1 ) ;
assign n76 =  ( n28 ) ? ( LB2D_shift_1 ) : ( n75 ) ;
assign n77 =  ( n23 ) ? ( LB2D_shift_0 ) : ( n76 ) ;
assign n78 =  ( n18 ) ? ( LB2D_shift_1 ) : ( n77 ) ;
assign n79 =  ( n9 ) ? ( LB2D_shift_1 ) : ( n78 ) ;
assign n80 =  ( n4 ) ? ( LB2D_shift_1 ) : ( n79 ) ;
assign n81 =  ( n31 ) ? ( LB2D_shift_2 ) : ( LB2D_shift_2 ) ;
assign n82 =  ( n28 ) ? ( LB2D_shift_2 ) : ( n81 ) ;
assign n83 =  ( n23 ) ? ( LB2D_shift_1 ) : ( n82 ) ;
assign n84 =  ( n18 ) ? ( LB2D_shift_2 ) : ( n83 ) ;
assign n85 =  ( n9 ) ? ( LB2D_shift_2 ) : ( n84 ) ;
assign n86 =  ( n4 ) ? ( LB2D_shift_2 ) : ( n85 ) ;
assign n87 =  ( n31 ) ? ( LB2D_shift_3 ) : ( LB2D_shift_3 ) ;
assign n88 =  ( n28 ) ? ( LB2D_shift_3 ) : ( n87 ) ;
assign n89 =  ( n23 ) ? ( LB2D_shift_2 ) : ( n88 ) ;
assign n90 =  ( n18 ) ? ( LB2D_shift_3 ) : ( n89 ) ;
assign n91 =  ( n9 ) ? ( LB2D_shift_3 ) : ( n90 ) ;
assign n92 =  ( n4 ) ? ( LB2D_shift_3 ) : ( n91 ) ;
assign n93 =  ( n31 ) ? ( LB2D_shift_4 ) : ( LB2D_shift_4 ) ;
assign n94 =  ( n28 ) ? ( LB2D_shift_4 ) : ( n93 ) ;
assign n95 =  ( n23 ) ? ( LB2D_shift_3 ) : ( n94 ) ;
assign n96 =  ( n18 ) ? ( LB2D_shift_4 ) : ( n95 ) ;
assign n97 =  ( n9 ) ? ( LB2D_shift_4 ) : ( n96 ) ;
assign n98 =  ( n4 ) ? ( LB2D_shift_4 ) : ( n97 ) ;
assign n99 =  ( n31 ) ? ( LB2D_shift_5 ) : ( LB2D_shift_5 ) ;
assign n100 =  ( n28 ) ? ( LB2D_shift_5 ) : ( n99 ) ;
assign n101 =  ( n23 ) ? ( LB2D_shift_4 ) : ( n100 ) ;
assign n102 =  ( n18 ) ? ( LB2D_shift_5 ) : ( n101 ) ;
assign n103 =  ( n9 ) ? ( LB2D_shift_5 ) : ( n102 ) ;
assign n104 =  ( n4 ) ? ( LB2D_shift_5 ) : ( n103 ) ;
assign n105 =  ( n31 ) ? ( LB2D_shift_6 ) : ( LB2D_shift_6 ) ;
assign n106 =  ( n28 ) ? ( LB2D_shift_6 ) : ( n105 ) ;
assign n107 =  ( n23 ) ? ( LB2D_shift_5 ) : ( n106 ) ;
assign n108 =  ( n18 ) ? ( LB2D_shift_6 ) : ( n107 ) ;
assign n109 =  ( n9 ) ? ( LB2D_shift_6 ) : ( n108 ) ;
assign n110 =  ( n4 ) ? ( LB2D_shift_6 ) : ( n109 ) ;
assign n111 =  ( n31 ) ? ( LB2D_shift_7 ) : ( LB2D_shift_7 ) ;
assign n112 =  ( n28 ) ? ( LB2D_shift_7 ) : ( n111 ) ;
assign n113 =  ( n23 ) ? ( LB2D_shift_6 ) : ( n112 ) ;
assign n114 =  ( n18 ) ? ( LB2D_shift_7 ) : ( n113 ) ;
assign n115 =  ( n9 ) ? ( LB2D_shift_7 ) : ( n114 ) ;
assign n116 =  ( n4 ) ? ( LB2D_shift_7 ) : ( n115 ) ;
assign n117 =  ( LB2D_shift_x ) < ( 9'd487 )  ;
assign n118 =  ( LB2D_shift_x ) + ( 9'd1 )  ;
assign n119 =  ( n117 ) ? ( n118 ) : ( 9'd0 ) ;
assign n120 =  ( n31 ) ? ( LB2D_shift_x ) : ( LB2D_shift_x ) ;
assign n121 =  ( n28 ) ? ( LB2D_shift_x ) : ( n120 ) ;
assign n122 =  ( n23 ) ? ( n119 ) : ( n121 ) ;
assign n123 =  ( n18 ) ? ( LB2D_shift_x ) : ( n122 ) ;
assign n124 =  ( n9 ) ? ( LB2D_shift_x ) : ( n123 ) ;
assign n125 =  ( n4 ) ? ( LB2D_shift_x ) : ( n124 ) ;
assign n126 =  ( LB2D_shift_y ) < ( 10'd487 )  ;
assign n127 =  ( LB2D_shift_y ) + ( 10'd1 )  ;
assign n128 =  ( n117 ) ? ( LB2D_shift_y ) : ( n127 ) ;
assign n129 =  ( n126 ) ? ( n128 ) : ( 10'd487 ) ;
assign n130 =  ( n31 ) ? ( LB2D_shift_y ) : ( LB2D_shift_y ) ;
assign n131 =  ( n28 ) ? ( LB2D_shift_y ) : ( n130 ) ;
assign n132 =  ( n23 ) ? ( n129 ) : ( n131 ) ;
assign n133 =  ( n18 ) ? ( LB2D_shift_y ) : ( n132 ) ;
assign n134 =  ( n9 ) ? ( LB2D_shift_y ) : ( n133 ) ;
assign n135 =  ( n4 ) ? ( LB2D_shift_y ) : ( n134 ) ;
assign n136 =  ( stencil_stream_full ) == ( 1'd1 )  ;
assign n137 =  ( n136 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_0 ) ;
assign n138 = gb_fun(n137) ;
assign n139 =  ( n31 ) ? ( arg_0_TDATA ) : ( arg_0_TDATA ) ;
assign n140 =  ( n28 ) ? ( arg_0_TDATA ) : ( n139 ) ;
assign n141 =  ( n23 ) ? ( arg_0_TDATA ) : ( n140 ) ;
assign n142 =  ( n18 ) ? ( n138 ) : ( n141 ) ;
assign n143 =  ( n9 ) ? ( arg_0_TDATA ) : ( n142 ) ;
assign n144 =  ( n4 ) ? ( arg_0_TDATA ) : ( n143 ) ;
assign n145 =  ( gb_pp_it_7 ) == ( 1'd1 )  ;
assign n146 =  ( n145 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n147 =  ( n31 ) ? ( arg_0_TVALID ) : ( arg_0_TVALID ) ;
assign n148 =  ( n28 ) ? ( arg_0_TVALID ) : ( n147 ) ;
assign n149 =  ( n23 ) ? ( arg_0_TVALID ) : ( n148 ) ;
assign n150 =  ( n18 ) ? ( n146 ) : ( n149 ) ;
assign n151 =  ( n9 ) ? ( arg_0_TVALID ) : ( n150 ) ;
assign n152 =  ( n4 ) ? ( 1'd0 ) : ( n151 ) ;
assign n153 =  ( n31 ) ? ( 1'd1 ) : ( arg_1_TREADY ) ;
assign n154 =  ( n28 ) ? ( arg_1_TREADY ) : ( n153 ) ;
assign n155 =  ( n23 ) ? ( arg_1_TREADY ) : ( n154 ) ;
assign n156 =  ( n18 ) ? ( arg_1_TREADY ) : ( n155 ) ;
assign n157 =  ( n9 ) ? ( 1'd0 ) : ( n156 ) ;
assign n158 =  ( n4 ) ? ( 1'd0 ) : ( n157 ) ;
assign n159 =  ( p_cnt ) + ( 19'd1 )  ;
assign n160 =  ( n159 ) == ( 19'd307200 )  ;
assign n161 =  ( n160 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n162 =  ( n18 ) ? ( n161 ) : ( gb_exit_it_1 ) ;
assign n163 =  ( n18 ) ? ( gb_exit_it_1 ) : ( gb_exit_it_2 ) ;
assign n164 =  ( n18 ) ? ( gb_exit_it_2 ) : ( gb_exit_it_3 ) ;
assign n165 =  ( n18 ) ? ( gb_exit_it_3 ) : ( gb_exit_it_4 ) ;
assign n166 =  ( n18 ) ? ( gb_exit_it_4 ) : ( gb_exit_it_5 ) ;
assign n167 =  ( n18 ) ? ( gb_exit_it_5 ) : ( gb_exit_it_6 ) ;
assign n168 =  ( n18 ) ? ( gb_exit_it_6 ) : ( gb_exit_it_7 ) ;
assign n169 =  ( n18 ) ? ( gb_exit_it_7 ) : ( gb_exit_it_8 ) ;
assign n170 =  ( n18 ) ? ( 1'd1 ) : ( gb_pp_it_1 ) ;
assign n171 =  ( n18 ) ? ( gb_pp_it_1 ) : ( gb_pp_it_2 ) ;
assign n172 =  ( n18 ) ? ( gb_pp_it_2 ) : ( gb_pp_it_3 ) ;
assign n173 =  ( n18 ) ? ( gb_pp_it_3 ) : ( gb_pp_it_4 ) ;
assign n174 =  ( n18 ) ? ( gb_pp_it_4 ) : ( gb_pp_it_5 ) ;
assign n175 =  ( n18 ) ? ( gb_pp_it_5 ) : ( gb_pp_it_6 ) ;
assign n176 =  ( n18 ) ? ( gb_pp_it_6 ) : ( gb_pp_it_7 ) ;
assign n177 =  ( n18 ) ? ( gb_pp_it_7 ) : ( gb_pp_it_8 ) ;
assign n178 =  ( n18 ) ? ( gb_pp_it_8 ) : ( gb_pp_it_9 ) ;
assign n179 =  ( n31 ) ? ( LB1D_buff ) : ( in_stream_buff_0 ) ;
assign n180 =  ( n28 ) ? ( in_stream_buff_0 ) : ( n179 ) ;
assign n181 =  ( n23 ) ? ( in_stream_buff_0 ) : ( n180 ) ;
assign n182 =  ( n18 ) ? ( in_stream_buff_0 ) : ( n181 ) ;
assign n183 =  ( n9 ) ? ( in_stream_buff_0 ) : ( n182 ) ;
assign n184 =  ( n4 ) ? ( in_stream_buff_0 ) : ( n183 ) ;
assign n185 =  ( n31 ) ? ( in_stream_buff_0 ) : ( in_stream_buff_1 ) ;
assign n186 =  ( n28 ) ? ( in_stream_buff_1 ) : ( n185 ) ;
assign n187 =  ( n23 ) ? ( in_stream_buff_1 ) : ( n186 ) ;
assign n188 =  ( n18 ) ? ( in_stream_buff_1 ) : ( n187 ) ;
assign n189 =  ( n9 ) ? ( in_stream_buff_1 ) : ( n188 ) ;
assign n190 =  ( n4 ) ? ( in_stream_buff_1 ) : ( n189 ) ;
assign n191 =  ( in_stream_full ) == ( 1'd1 )  ;
assign n192 =  ( n191 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n193 =  ( n31 ) ? ( 1'd0 ) : ( in_stream_empty ) ;
assign n194 =  ( n28 ) ? ( n192 ) : ( n193 ) ;
assign n195 =  ( n23 ) ? ( in_stream_empty ) : ( n194 ) ;
assign n196 =  ( n18 ) ? ( in_stream_empty ) : ( n195 ) ;
assign n197 =  ( n9 ) ? ( in_stream_empty ) : ( n196 ) ;
assign n198 =  ( n4 ) ? ( in_stream_empty ) : ( n197 ) ;
assign n199 =  ( in_stream_empty ) == ( 1'd1 )  ;
assign n200 =  ( n199 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n201 =  ( n31 ) ? ( n200 ) : ( in_stream_full ) ;
assign n202 =  ( n28 ) ? ( 1'd0 ) : ( n201 ) ;
assign n203 =  ( n23 ) ? ( in_stream_full ) : ( n202 ) ;
assign n204 =  ( n18 ) ? ( in_stream_full ) : ( n203 ) ;
assign n205 =  ( n9 ) ? ( in_stream_full ) : ( n204 ) ;
assign n206 =  ( n4 ) ? ( in_stream_full ) : ( n205 ) ;
assign n207 =  ( p_cnt ) < ( 19'd307200 )  ;
assign n208 =  ( n207 ) ? ( n159 ) : ( 19'd307200 ) ;
assign n209 =  ( n18 ) ? ( n208 ) : ( p_cnt ) ;
assign n210 =  ( n191 ) ? ( in_stream_buff_1 ) : ( in_stream_buff_0 ) ;
assign n211 =  ( LB2D_proc_w ) == ( 64'd0 )  ;
assign n212 =  (  LB2D_proc_7 [ LB2D_proc_x ] )  ;
assign n213 =  ( LB2D_proc_w ) == ( 64'd1 )  ;
assign n214 =  (  LB2D_proc_0 [ LB2D_proc_x ] )  ;
assign n215 =  ( LB2D_proc_w ) == ( 64'd2 )  ;
assign n216 =  (  LB2D_proc_1 [ LB2D_proc_x ] )  ;
assign n217 =  ( LB2D_proc_w ) == ( 64'd3 )  ;
assign n218 =  (  LB2D_proc_2 [ LB2D_proc_x ] )  ;
assign n219 =  ( LB2D_proc_w ) == ( 64'd4 )  ;
assign n220 =  (  LB2D_proc_3 [ LB2D_proc_x ] )  ;
assign n221 =  ( LB2D_proc_w ) == ( 64'd5 )  ;
assign n222 =  (  LB2D_proc_4 [ LB2D_proc_x ] )  ;
assign n223 =  ( LB2D_proc_w ) == ( 64'd6 )  ;
assign n224 =  (  LB2D_proc_5 [ LB2D_proc_x ] )  ;
assign n225 =  (  LB2D_proc_6 [ LB2D_proc_x ] )  ;
assign n226 =  ( n223 ) ? ( n224 ) : ( n225 ) ;
assign n227 =  ( n221 ) ? ( n222 ) : ( n226 ) ;
assign n228 =  ( n219 ) ? ( n220 ) : ( n227 ) ;
assign n229 =  ( n217 ) ? ( n218 ) : ( n228 ) ;
assign n230 =  ( n215 ) ? ( n216 ) : ( n229 ) ;
assign n231 =  ( n213 ) ? ( n214 ) : ( n230 ) ;
assign n232 =  ( n211 ) ? ( n212 ) : ( n231 ) ;
assign n233 =  ( n223 ) ? ( n222 ) : ( n224 ) ;
assign n234 =  ( n221 ) ? ( n220 ) : ( n233 ) ;
assign n235 =  ( n219 ) ? ( n218 ) : ( n234 ) ;
assign n236 =  ( n217 ) ? ( n216 ) : ( n235 ) ;
assign n237 =  ( n215 ) ? ( n214 ) : ( n236 ) ;
assign n238 =  ( n213 ) ? ( n212 ) : ( n237 ) ;
assign n239 =  ( n211 ) ? ( n225 ) : ( n238 ) ;
assign n240 =  ( n223 ) ? ( n220 ) : ( n222 ) ;
assign n241 =  ( n221 ) ? ( n218 ) : ( n240 ) ;
assign n242 =  ( n219 ) ? ( n216 ) : ( n241 ) ;
assign n243 =  ( n217 ) ? ( n214 ) : ( n242 ) ;
assign n244 =  ( n215 ) ? ( n212 ) : ( n243 ) ;
assign n245 =  ( n213 ) ? ( n225 ) : ( n244 ) ;
assign n246 =  ( n211 ) ? ( n224 ) : ( n245 ) ;
assign n247 =  ( n223 ) ? ( n218 ) : ( n220 ) ;
assign n248 =  ( n221 ) ? ( n216 ) : ( n247 ) ;
assign n249 =  ( n219 ) ? ( n214 ) : ( n248 ) ;
assign n250 =  ( n217 ) ? ( n212 ) : ( n249 ) ;
assign n251 =  ( n215 ) ? ( n225 ) : ( n250 ) ;
assign n252 =  ( n213 ) ? ( n224 ) : ( n251 ) ;
assign n253 =  ( n211 ) ? ( n222 ) : ( n252 ) ;
assign n254 =  ( n223 ) ? ( n216 ) : ( n218 ) ;
assign n255 =  ( n221 ) ? ( n214 ) : ( n254 ) ;
assign n256 =  ( n219 ) ? ( n212 ) : ( n255 ) ;
assign n257 =  ( n217 ) ? ( n225 ) : ( n256 ) ;
assign n258 =  ( n215 ) ? ( n224 ) : ( n257 ) ;
assign n259 =  ( n213 ) ? ( n222 ) : ( n258 ) ;
assign n260 =  ( n211 ) ? ( n220 ) : ( n259 ) ;
assign n261 =  ( n223 ) ? ( n214 ) : ( n216 ) ;
assign n262 =  ( n221 ) ? ( n212 ) : ( n261 ) ;
assign n263 =  ( n219 ) ? ( n225 ) : ( n262 ) ;
assign n264 =  ( n217 ) ? ( n224 ) : ( n263 ) ;
assign n265 =  ( n215 ) ? ( n222 ) : ( n264 ) ;
assign n266 =  ( n213 ) ? ( n220 ) : ( n265 ) ;
assign n267 =  ( n211 ) ? ( n218 ) : ( n266 ) ;
assign n268 =  ( n223 ) ? ( n212 ) : ( n214 ) ;
assign n269 =  ( n221 ) ? ( n225 ) : ( n268 ) ;
assign n270 =  ( n219 ) ? ( n224 ) : ( n269 ) ;
assign n271 =  ( n217 ) ? ( n222 ) : ( n270 ) ;
assign n272 =  ( n215 ) ? ( n220 ) : ( n271 ) ;
assign n273 =  ( n213 ) ? ( n218 ) : ( n272 ) ;
assign n274 =  ( n211 ) ? ( n216 ) : ( n273 ) ;
assign n275 =  ( n223 ) ? ( n225 ) : ( n212 ) ;
assign n276 =  ( n221 ) ? ( n224 ) : ( n275 ) ;
assign n277 =  ( n219 ) ? ( n222 ) : ( n276 ) ;
assign n278 =  ( n217 ) ? ( n220 ) : ( n277 ) ;
assign n279 =  ( n215 ) ? ( n218 ) : ( n278 ) ;
assign n280 =  ( n213 ) ? ( n216 ) : ( n279 ) ;
assign n281 =  ( n211 ) ? ( n214 ) : ( n280 ) ;
assign n282 =  { ( n274 ) , ( n281 ) }  ;
assign n283 =  { ( n267 ) , ( n282 ) }  ;
assign n284 =  { ( n260 ) , ( n283 ) }  ;
assign n285 =  { ( n253 ) , ( n284 ) }  ;
assign n286 =  { ( n246 ) , ( n285 ) }  ;
assign n287 =  { ( n239 ) , ( n286 ) }  ;
assign n288 =  { ( n232 ) , ( n287 ) }  ;
assign n289 =  { ( n210 ) , ( n288 ) }  ;
assign n290 =  ( n26 ) ? ( slice_stream_buff_0 ) : ( n289 ) ;
assign n291 =  ( n31 ) ? ( slice_stream_buff_0 ) : ( slice_stream_buff_0 ) ;
assign n292 =  ( n28 ) ? ( n290 ) : ( n291 ) ;
assign n293 =  ( n23 ) ? ( slice_stream_buff_0 ) : ( n292 ) ;
assign n294 =  ( n18 ) ? ( slice_stream_buff_0 ) : ( n293 ) ;
assign n295 =  ( n9 ) ? ( slice_stream_buff_0 ) : ( n294 ) ;
assign n296 =  ( n4 ) ? ( slice_stream_buff_0 ) : ( n295 ) ;
assign n297 =  ( n26 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n298 =  ( n31 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_1 ) ;
assign n299 =  ( n28 ) ? ( n297 ) : ( n298 ) ;
assign n300 =  ( n23 ) ? ( slice_stream_buff_1 ) : ( n299 ) ;
assign n301 =  ( n18 ) ? ( slice_stream_buff_1 ) : ( n300 ) ;
assign n302 =  ( n9 ) ? ( slice_stream_buff_1 ) : ( n301 ) ;
assign n303 =  ( n4 ) ? ( slice_stream_buff_1 ) : ( n302 ) ;
assign n304 =  ( n67 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n305 =  ( n26 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n306 =  ( n31 ) ? ( slice_stream_empty ) : ( slice_stream_empty ) ;
assign n307 =  ( n28 ) ? ( n305 ) : ( n306 ) ;
assign n308 =  ( n23 ) ? ( n304 ) : ( n307 ) ;
assign n309 =  ( n18 ) ? ( slice_stream_empty ) : ( n308 ) ;
assign n310 =  ( n9 ) ? ( slice_stream_empty ) : ( n309 ) ;
assign n311 =  ( n4 ) ? ( slice_stream_empty ) : ( n310 ) ;
assign n312 =  ( slice_stream_empty ) == ( 1'd1 )  ;
assign n313 =  ( n312 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n314 =  ( n26 ) ? ( 1'd0 ) : ( n313 ) ;
assign n315 =  ( n31 ) ? ( slice_stream_full ) : ( slice_stream_full ) ;
assign n316 =  ( n28 ) ? ( n314 ) : ( n315 ) ;
assign n317 =  ( n23 ) ? ( 1'd0 ) : ( n316 ) ;
assign n318 =  ( n18 ) ? ( slice_stream_full ) : ( n317 ) ;
assign n319 =  ( n9 ) ? ( slice_stream_full ) : ( n318 ) ;
assign n320 =  ( n4 ) ? ( slice_stream_full ) : ( n319 ) ;
assign n321 =  ( LB2D_shift_x ) >= ( 9'd8 )  ;
assign n322 = n68[71:64] ;
assign n323 = LB2D_shift_0[71:64] ;
assign n324 = LB2D_shift_1[71:64] ;
assign n325 = LB2D_shift_2[71:64] ;
assign n326 = LB2D_shift_3[71:64] ;
assign n327 = LB2D_shift_4[71:64] ;
assign n328 = LB2D_shift_5[71:64] ;
assign n329 = LB2D_shift_6[71:64] ;
assign n330 = LB2D_shift_7[71:64] ;
assign n331 =  { ( n329 ) , ( n330 ) }  ;
assign n332 =  { ( n328 ) , ( n331 ) }  ;
assign n333 =  { ( n327 ) , ( n332 ) }  ;
assign n334 =  { ( n326 ) , ( n333 ) }  ;
assign n335 =  { ( n325 ) , ( n334 ) }  ;
assign n336 =  { ( n324 ) , ( n335 ) }  ;
assign n337 =  { ( n323 ) , ( n336 ) }  ;
assign n338 =  { ( n322 ) , ( n337 ) }  ;
assign n339 = n68[63:56] ;
assign n340 = LB2D_shift_0[63:56] ;
assign n341 = LB2D_shift_1[63:56] ;
assign n342 = LB2D_shift_2[63:56] ;
assign n343 = LB2D_shift_3[63:56] ;
assign n344 = LB2D_shift_4[63:56] ;
assign n345 = LB2D_shift_5[63:56] ;
assign n346 = LB2D_shift_6[63:56] ;
assign n347 = LB2D_shift_7[63:56] ;
assign n348 =  { ( n346 ) , ( n347 ) }  ;
assign n349 =  { ( n345 ) , ( n348 ) }  ;
assign n350 =  { ( n344 ) , ( n349 ) }  ;
assign n351 =  { ( n343 ) , ( n350 ) }  ;
assign n352 =  { ( n342 ) , ( n351 ) }  ;
assign n353 =  { ( n341 ) , ( n352 ) }  ;
assign n354 =  { ( n340 ) , ( n353 ) }  ;
assign n355 =  { ( n339 ) , ( n354 ) }  ;
assign n356 = n68[55:48] ;
assign n357 = LB2D_shift_0[55:48] ;
assign n358 = LB2D_shift_1[55:48] ;
assign n359 = LB2D_shift_2[55:48] ;
assign n360 = LB2D_shift_3[55:48] ;
assign n361 = LB2D_shift_4[55:48] ;
assign n362 = LB2D_shift_5[55:48] ;
assign n363 = LB2D_shift_6[55:48] ;
assign n364 = LB2D_shift_7[55:48] ;
assign n365 =  { ( n363 ) , ( n364 ) }  ;
assign n366 =  { ( n362 ) , ( n365 ) }  ;
assign n367 =  { ( n361 ) , ( n366 ) }  ;
assign n368 =  { ( n360 ) , ( n367 ) }  ;
assign n369 =  { ( n359 ) , ( n368 ) }  ;
assign n370 =  { ( n358 ) , ( n369 ) }  ;
assign n371 =  { ( n357 ) , ( n370 ) }  ;
assign n372 =  { ( n356 ) , ( n371 ) }  ;
assign n373 = n68[47:40] ;
assign n374 = LB2D_shift_0[47:40] ;
assign n375 = LB2D_shift_1[47:40] ;
assign n376 = LB2D_shift_2[47:40] ;
assign n377 = LB2D_shift_3[47:40] ;
assign n378 = LB2D_shift_4[47:40] ;
assign n379 = LB2D_shift_5[47:40] ;
assign n380 = LB2D_shift_6[47:40] ;
assign n381 = LB2D_shift_7[47:40] ;
assign n382 =  { ( n380 ) , ( n381 ) }  ;
assign n383 =  { ( n379 ) , ( n382 ) }  ;
assign n384 =  { ( n378 ) , ( n383 ) }  ;
assign n385 =  { ( n377 ) , ( n384 ) }  ;
assign n386 =  { ( n376 ) , ( n385 ) }  ;
assign n387 =  { ( n375 ) , ( n386 ) }  ;
assign n388 =  { ( n374 ) , ( n387 ) }  ;
assign n389 =  { ( n373 ) , ( n388 ) }  ;
assign n390 = n68[39:32] ;
assign n391 = LB2D_shift_0[39:32] ;
assign n392 = LB2D_shift_1[39:32] ;
assign n393 = LB2D_shift_2[39:32] ;
assign n394 = LB2D_shift_3[39:32] ;
assign n395 = LB2D_shift_4[39:32] ;
assign n396 = LB2D_shift_5[39:32] ;
assign n397 = LB2D_shift_6[39:32] ;
assign n398 = LB2D_shift_7[39:32] ;
assign n399 =  { ( n397 ) , ( n398 ) }  ;
assign n400 =  { ( n396 ) , ( n399 ) }  ;
assign n401 =  { ( n395 ) , ( n400 ) }  ;
assign n402 =  { ( n394 ) , ( n401 ) }  ;
assign n403 =  { ( n393 ) , ( n402 ) }  ;
assign n404 =  { ( n392 ) , ( n403 ) }  ;
assign n405 =  { ( n391 ) , ( n404 ) }  ;
assign n406 =  { ( n390 ) , ( n405 ) }  ;
assign n407 = n68[31:24] ;
assign n408 = LB2D_shift_0[31:24] ;
assign n409 = LB2D_shift_1[31:24] ;
assign n410 = LB2D_shift_2[31:24] ;
assign n411 = LB2D_shift_3[31:24] ;
assign n412 = LB2D_shift_4[31:24] ;
assign n413 = LB2D_shift_5[31:24] ;
assign n414 = LB2D_shift_6[31:24] ;
assign n415 = LB2D_shift_7[31:24] ;
assign n416 =  { ( n414 ) , ( n415 ) }  ;
assign n417 =  { ( n413 ) , ( n416 ) }  ;
assign n418 =  { ( n412 ) , ( n417 ) }  ;
assign n419 =  { ( n411 ) , ( n418 ) }  ;
assign n420 =  { ( n410 ) , ( n419 ) }  ;
assign n421 =  { ( n409 ) , ( n420 ) }  ;
assign n422 =  { ( n408 ) , ( n421 ) }  ;
assign n423 =  { ( n407 ) , ( n422 ) }  ;
assign n424 = n68[23:16] ;
assign n425 = LB2D_shift_0[23:16] ;
assign n426 = LB2D_shift_1[23:16] ;
assign n427 = LB2D_shift_2[23:16] ;
assign n428 = LB2D_shift_3[23:16] ;
assign n429 = LB2D_shift_4[23:16] ;
assign n430 = LB2D_shift_5[23:16] ;
assign n431 = LB2D_shift_6[23:16] ;
assign n432 = LB2D_shift_7[23:16] ;
assign n433 =  { ( n431 ) , ( n432 ) }  ;
assign n434 =  { ( n430 ) , ( n433 ) }  ;
assign n435 =  { ( n429 ) , ( n434 ) }  ;
assign n436 =  { ( n428 ) , ( n435 ) }  ;
assign n437 =  { ( n427 ) , ( n436 ) }  ;
assign n438 =  { ( n426 ) , ( n437 ) }  ;
assign n439 =  { ( n425 ) , ( n438 ) }  ;
assign n440 =  { ( n424 ) , ( n439 ) }  ;
assign n441 = n68[15:8] ;
assign n442 = LB2D_shift_0[15:8] ;
assign n443 = LB2D_shift_1[15:8] ;
assign n444 = LB2D_shift_2[15:8] ;
assign n445 = LB2D_shift_3[15:8] ;
assign n446 = LB2D_shift_4[15:8] ;
assign n447 = LB2D_shift_5[15:8] ;
assign n448 = LB2D_shift_6[15:8] ;
assign n449 = LB2D_shift_7[15:8] ;
assign n450 =  { ( n448 ) , ( n449 ) }  ;
assign n451 =  { ( n447 ) , ( n450 ) }  ;
assign n452 =  { ( n446 ) , ( n451 ) }  ;
assign n453 =  { ( n445 ) , ( n452 ) }  ;
assign n454 =  { ( n444 ) , ( n453 ) }  ;
assign n455 =  { ( n443 ) , ( n454 ) }  ;
assign n456 =  { ( n442 ) , ( n455 ) }  ;
assign n457 =  { ( n441 ) , ( n456 ) }  ;
assign n458 = n68[7:0] ;
assign n459 = LB2D_shift_0[7:0] ;
assign n460 = LB2D_shift_1[7:0] ;
assign n461 = LB2D_shift_2[7:0] ;
assign n462 = LB2D_shift_3[7:0] ;
assign n463 = LB2D_shift_4[7:0] ;
assign n464 = LB2D_shift_5[7:0] ;
assign n465 = LB2D_shift_6[7:0] ;
assign n466 = LB2D_shift_7[7:0] ;
assign n467 =  { ( n465 ) , ( n466 ) }  ;
assign n468 =  { ( n464 ) , ( n467 ) }  ;
assign n469 =  { ( n463 ) , ( n468 ) }  ;
assign n470 =  { ( n462 ) , ( n469 ) }  ;
assign n471 =  { ( n461 ) , ( n470 ) }  ;
assign n472 =  { ( n460 ) , ( n471 ) }  ;
assign n473 =  { ( n459 ) , ( n472 ) }  ;
assign n474 =  { ( n458 ) , ( n473 ) }  ;
assign n475 =  { ( n457 ) , ( n474 ) }  ;
assign n476 =  { ( n440 ) , ( n475 ) }  ;
assign n477 =  { ( n423 ) , ( n476 ) }  ;
assign n478 =  { ( n406 ) , ( n477 ) }  ;
assign n479 =  { ( n389 ) , ( n478 ) }  ;
assign n480 =  { ( n372 ) , ( n479 ) }  ;
assign n481 =  { ( n355 ) , ( n480 ) }  ;
assign n482 =  { ( n338 ) , ( n481 ) }  ;
assign n483 =  ( n321 ) ? ( n482 ) : ( stencil_stream_buff_0 ) ;
assign n484 =  ( n31 ) ? ( stencil_stream_buff_0 ) : ( stencil_stream_buff_0 ) ;
assign n485 =  ( n28 ) ? ( stencil_stream_buff_0 ) : ( n484 ) ;
assign n486 =  ( n23 ) ? ( n483 ) : ( n485 ) ;
assign n487 =  ( n18 ) ? ( stencil_stream_buff_0 ) : ( n486 ) ;
assign n488 =  ( n9 ) ? ( stencil_stream_buff_0 ) : ( n487 ) ;
assign n489 =  ( n4 ) ? ( stencil_stream_buff_0 ) : ( n488 ) ;
assign n490 =  ( n31 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_1 ) ;
assign n491 =  ( n28 ) ? ( stencil_stream_buff_1 ) : ( n490 ) ;
assign n492 =  ( n23 ) ? ( stencil_stream_buff_0 ) : ( n491 ) ;
assign n493 =  ( n18 ) ? ( stencil_stream_buff_1 ) : ( n492 ) ;
assign n494 =  ( n9 ) ? ( stencil_stream_buff_1 ) : ( n493 ) ;
assign n495 =  ( n4 ) ? ( stencil_stream_buff_1 ) : ( n494 ) ;
assign n496 =  ( n136 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n497 =  ( n21 ) ? ( stencil_stream_empty ) : ( 1'd0 ) ;
assign n498 =  ( n31 ) ? ( stencil_stream_empty ) : ( stencil_stream_empty ) ;
assign n499 =  ( n28 ) ? ( stencil_stream_empty ) : ( n498 ) ;
assign n500 =  ( n23 ) ? ( n497 ) : ( n499 ) ;
assign n501 =  ( n18 ) ? ( n496 ) : ( n500 ) ;
assign n502 =  ( n9 ) ? ( stencil_stream_empty ) : ( n501 ) ;
assign n503 =  ( n4 ) ? ( stencil_stream_empty ) : ( n502 ) ;
assign n504 =  ( n14 ) ? ( 1'd0 ) : ( 1'd0 ) ;
assign n505 =  ( stencil_stream_empty ) == ( 1'd1 )  ;
assign n506 =  ( n505 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n507 =  ( n21 ) ? ( stencil_stream_full ) : ( n506 ) ;
assign n508 =  ( n31 ) ? ( stencil_stream_full ) : ( stencil_stream_full ) ;
assign n509 =  ( n28 ) ? ( stencil_stream_full ) : ( n508 ) ;
assign n510 =  ( n23 ) ? ( n507 ) : ( n509 ) ;
assign n511 =  ( n18 ) ? ( n504 ) : ( n510 ) ;
assign n512 =  ( n9 ) ? ( stencil_stream_full ) : ( n511 ) ;
assign n513 =  ( n4 ) ? ( stencil_stream_full ) : ( n512 ) ;
assign n514 = ~ ( n4 ) ;
assign n515 = ~ ( n9 ) ;
assign n516 =  ( n514 ) & ( n515 )  ;
assign n517 = ~ ( n18 ) ;
assign n518 =  ( n516 ) & ( n517 )  ;
assign n519 = ~ ( n23 ) ;
assign n520 =  ( n518 ) & ( n519 )  ;
assign n521 = ~ ( n28 ) ;
assign n522 =  ( n520 ) & ( n521 )  ;
assign n523 = ~ ( n31 ) ;
assign n524 =  ( n522 ) & ( n523 )  ;
assign n525 =  ( n522 ) & ( n31 )  ;
assign n526 =  ( n520 ) & ( n28 )  ;
assign n527 = ~ ( n211 ) ;
assign n528 =  ( n526 ) & ( n527 )  ;
assign n529 =  ( n526 ) & ( n211 )  ;
assign n530 =  ( n518 ) & ( n23 )  ;
assign n531 =  ( n516 ) & ( n18 )  ;
assign n532 =  ( n514 ) & ( n9 )  ;
assign LB2D_proc_0_addr0 = n529 ? (LB2D_proc_x) : (0);
assign LB2D_proc_0_data0 = n529 ? (n210) : (LB2D_proc_0[0]);
assign n533 = ~ ( n213 ) ;
assign n534 =  ( n526 ) & ( n533 )  ;
assign n535 =  ( n526 ) & ( n213 )  ;
assign LB2D_proc_1_addr0 = n535 ? (LB2D_proc_x) : (0);
assign LB2D_proc_1_data0 = n535 ? (n210) : (LB2D_proc_1[0]);
assign n536 = ~ ( n215 ) ;
assign n537 =  ( n526 ) & ( n536 )  ;
assign n538 =  ( n526 ) & ( n215 )  ;
assign LB2D_proc_2_addr0 = n538 ? (LB2D_proc_x) : (0);
assign LB2D_proc_2_data0 = n538 ? (n210) : (LB2D_proc_2[0]);
assign n539 = ~ ( n217 ) ;
assign n540 =  ( n526 ) & ( n539 )  ;
assign n541 =  ( n526 ) & ( n217 )  ;
assign LB2D_proc_3_addr0 = n541 ? (LB2D_proc_x) : (0);
assign LB2D_proc_3_data0 = n541 ? (n210) : (LB2D_proc_3[0]);
assign n542 = ~ ( n219 ) ;
assign n543 =  ( n526 ) & ( n542 )  ;
assign n544 =  ( n526 ) & ( n219 )  ;
assign LB2D_proc_4_addr0 = n544 ? (LB2D_proc_x) : (0);
assign LB2D_proc_4_data0 = n544 ? (n210) : (LB2D_proc_4[0]);
assign n545 = ~ ( n221 ) ;
assign n546 =  ( n526 ) & ( n545 )  ;
assign n547 =  ( n526 ) & ( n221 )  ;
assign LB2D_proc_5_addr0 = n547 ? (LB2D_proc_x) : (0);
assign LB2D_proc_5_data0 = n547 ? (n210) : (LB2D_proc_5[0]);
assign n548 = ~ ( n223 ) ;
assign n549 =  ( n526 ) & ( n548 )  ;
assign n550 =  ( n526 ) & ( n223 )  ;
assign LB2D_proc_6_addr0 = n550 ? (LB2D_proc_x) : (0);
assign LB2D_proc_6_data0 = n550 ? (n210) : (LB2D_proc_6[0]);
assign n551 =  ( LB2D_proc_w ) == ( 64'd7 )  ;
assign n552 = ~ ( n551 ) ;
assign n553 =  ( n526 ) & ( n552 )  ;
assign n554 =  ( n526 ) & ( n551 )  ;
assign LB2D_proc_7_addr0 = n554 ? (LB2D_proc_x) : (0);
assign LB2D_proc_7_data0 = n554 ? (n210) : (LB2D_proc_7[0]);
function [7:0] gb_fun ;
input [647:0] arg0;
    begin
//TODO: Add the specific function HERE.    end
endfunction

always @(posedge clk) begin
   if(rst) begin
       LB1D_buff <= LB1D_buff;
       LB2D_proc_w <= LB2D_proc_w;
       LB2D_proc_x <= LB2D_proc_x;
       LB2D_proc_y <= LB2D_proc_y;
       LB2D_shift_0 <= LB2D_shift_0;
       LB2D_shift_1 <= LB2D_shift_1;
       LB2D_shift_2 <= LB2D_shift_2;
       LB2D_shift_3 <= LB2D_shift_3;
       LB2D_shift_4 <= LB2D_shift_4;
       LB2D_shift_5 <= LB2D_shift_5;
       LB2D_shift_6 <= LB2D_shift_6;
       LB2D_shift_7 <= LB2D_shift_7;
       LB2D_shift_x <= LB2D_shift_x;
       LB2D_shift_y <= LB2D_shift_y;
       arg_0_TDATA <= arg_0_TDATA;
       arg_0_TVALID <= arg_0_TVALID;
       arg_1_TREADY <= arg_1_TREADY;
       gb_exit_it_1 <= gb_exit_it_1;
       gb_exit_it_2 <= gb_exit_it_2;
       gb_exit_it_3 <= gb_exit_it_3;
       gb_exit_it_4 <= gb_exit_it_4;
       gb_exit_it_5 <= gb_exit_it_5;
       gb_exit_it_6 <= gb_exit_it_6;
       gb_exit_it_7 <= gb_exit_it_7;
       gb_exit_it_8 <= gb_exit_it_8;
       gb_pp_it_1 <= gb_pp_it_1;
       gb_pp_it_2 <= gb_pp_it_2;
       gb_pp_it_3 <= gb_pp_it_3;
       gb_pp_it_4 <= gb_pp_it_4;
       gb_pp_it_5 <= gb_pp_it_5;
       gb_pp_it_6 <= gb_pp_it_6;
       gb_pp_it_7 <= gb_pp_it_7;
       gb_pp_it_8 <= gb_pp_it_8;
       gb_pp_it_9 <= gb_pp_it_9;
       in_stream_buff_0 <= in_stream_buff_0;
       in_stream_buff_1 <= in_stream_buff_1;
       in_stream_empty <= in_stream_empty;
       in_stream_full <= in_stream_full;
       p_cnt <= p_cnt;
       slice_stream_buff_0 <= slice_stream_buff_0;
       slice_stream_buff_1 <= slice_stream_buff_1;
       slice_stream_empty <= slice_stream_empty;
       slice_stream_full <= slice_stream_full;
       stencil_stream_buff_0 <= stencil_stream_buff_0;
       stencil_stream_buff_1 <= stencil_stream_buff_1;
       stencil_stream_empty <= stencil_stream_empty;
       stencil_stream_full <= stencil_stream_full;
   end
   else if(step) begin
       LB1D_buff <= n37;
       LB2D_proc_w <= n48;
       LB2D_proc_x <= n56;
       LB2D_proc_y <= n66;
       LB2D_shift_0 <= n74;
       LB2D_shift_1 <= n80;
       LB2D_shift_2 <= n86;
       LB2D_shift_3 <= n92;
       LB2D_shift_4 <= n98;
       LB2D_shift_5 <= n104;
       LB2D_shift_6 <= n110;
       LB2D_shift_7 <= n116;
       LB2D_shift_x <= n125;
       LB2D_shift_y <= n135;
       arg_0_TDATA <= n144;
       arg_0_TVALID <= n152;
       arg_1_TREADY <= n158;
       gb_exit_it_1 <= n162;
       gb_exit_it_2 <= n163;
       gb_exit_it_3 <= n164;
       gb_exit_it_4 <= n165;
       gb_exit_it_5 <= n166;
       gb_exit_it_6 <= n167;
       gb_exit_it_7 <= n168;
       gb_exit_it_8 <= n169;
       gb_pp_it_1 <= n170;
       gb_pp_it_2 <= n171;
       gb_pp_it_3 <= n172;
       gb_pp_it_4 <= n173;
       gb_pp_it_5 <= n174;
       gb_pp_it_6 <= n175;
       gb_pp_it_7 <= n176;
       gb_pp_it_8 <= n177;
       gb_pp_it_9 <= n178;
       in_stream_buff_0 <= n184;
       in_stream_buff_1 <= n190;
       in_stream_empty <= n198;
       in_stream_full <= n206;
       p_cnt <= n209;
       slice_stream_buff_0 <= n296;
       slice_stream_buff_1 <= n303;
       slice_stream_empty <= n311;
       slice_stream_full <= n320;
       stencil_stream_buff_0 <= n489;
       stencil_stream_buff_1 <= n495;
       stencil_stream_empty <= n503;
       stencil_stream_full <= n513;
       LB2D_proc_0 [ LB2D_proc_0_addr0 ] <= LB2D_proc_0_data0;
       LB2D_proc_1 [ LB2D_proc_1_addr0 ] <= LB2D_proc_1_data0;
       LB2D_proc_2 [ LB2D_proc_2_addr0 ] <= LB2D_proc_2_data0;
       LB2D_proc_3 [ LB2D_proc_3_addr0 ] <= LB2D_proc_3_data0;
       LB2D_proc_4 [ LB2D_proc_4_addr0 ] <= LB2D_proc_4_data0;
       LB2D_proc_5 [ LB2D_proc_5_addr0 ] <= LB2D_proc_5_data0;
       LB2D_proc_6 [ LB2D_proc_6_addr0 ] <= LB2D_proc_6_data0;
       LB2D_proc_7 [ LB2D_proc_7_addr0 ] <= LB2D_proc_7_data0;
   end
end
endmodule
