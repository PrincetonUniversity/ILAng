module SPEC_A(
arg_0_TREADY,
arg_1_TDATA,
arg_1_TVALID,
RAM_w,
RAM_x,
RAM_y,
arg_0_TDATA,
arg_0_TVALID,
arg_1_TREADY,
cur_pix,
gbit,
pre_pix,
proc_in,
st_ready,
stencil_0,
stencil_1,
stencil_2,
stencil_3,
stencil_4,
stencil_5,
stencil_6,
stencil_7,
stencil_8,
clk,rst,
step
);
input            arg_0_TREADY;
input      [7:0] arg_1_TDATA;
input            arg_1_TVALID;
input clk;
input rst;
input step;
output      [2:0] RAM_w;
output      [8:0] RAM_x;
output      [9:0] RAM_y;
output      [7:0] arg_0_TDATA;
output            arg_0_TVALID;
output            arg_1_TREADY;
output      [7:0] cur_pix;
output      [3:0] gbit;
output      [7:0] pre_pix;
output    [647:0] proc_in;
output            st_ready;
output     [71:0] stencil_0;
output     [71:0] stencil_1;
output     [71:0] stencil_2;
output     [71:0] stencil_3;
output     [71:0] stencil_4;
output     [71:0] stencil_5;
output     [71:0] stencil_6;
output     [71:0] stencil_7;
output     [71:0] stencil_8;
reg      [2:0] RAM_w;
reg      [8:0] RAM_x;
reg      [9:0] RAM_y;
reg      [7:0] arg_0_TDATA;
reg            arg_0_TVALID;
reg            arg_1_TREADY;
reg      [7:0] cur_pix;
reg      [3:0] gbit;
reg      [7:0] pre_pix;
reg    [647:0] proc_in;
reg            st_ready;
reg     [71:0] stencil_0;
reg     [71:0] stencil_1;
reg     [71:0] stencil_2;
reg     [71:0] stencil_3;
reg     [71:0] stencil_4;
reg     [71:0] stencil_5;
reg     [71:0] stencil_6;
reg     [71:0] stencil_7;
reg     [71:0] stencil_8;
wire            arg_0_TREADY;
wire      [7:0] arg_1_TDATA;
wire            arg_1_TVALID;
wire            n0;
wire            n1;
wire            n2;
wire            n3;
wire            n4;
wire            n5;
wire            n6;
wire            n7;
wire            n8;
wire            n9;
wire            n10;
wire            n11;
wire            n12;
wire            n13;
wire            n14;
wire            n15;
wire            n16;
wire            n17;
wire            n18;
wire            n19;
wire            n20;
wire      [2:0] n21;
wire      [2:0] n22;
wire      [2:0] n23;
wire            n24;
wire            n25;
wire            n26;
wire            n27;
wire            n28;
wire            n29;
wire      [2:0] n30;
wire      [2:0] n31;
wire      [2:0] n32;
wire      [2:0] n33;
wire      [2:0] n34;
wire      [8:0] n35;
wire      [8:0] n36;
wire      [8:0] n37;
wire      [8:0] n38;
wire      [8:0] n39;
wire      [8:0] n40;
wire      [8:0] n41;
wire            n42;
wire      [9:0] n43;
wire      [9:0] n44;
wire      [9:0] n45;
wire      [9:0] n46;
wire      [9:0] n47;
wire      [9:0] n48;
wire      [9:0] n49;
wire      [9:0] n50;
wire            n51;
wire            n52;
wire            n53;
wire            n54;
wire            n55;
wire            n56;
wire            n57;
wire            n58;
wire      [7:0] n59;
wire      [7:0] n60;
wire      [7:0] n61;
wire      [7:0] n62;
wire      [7:0] n63;
wire      [7:0] n64;
wire      [7:0] n65;
wire      [7:0] n66;
wire      [7:0] n67;
wire     [15:0] n68;
wire     [23:0] n69;
wire     [31:0] n70;
wire     [39:0] n71;
wire     [47:0] n72;
wire     [55:0] n73;
wire     [63:0] n74;
wire     [71:0] n75;
wire      [7:0] n76;
wire      [7:0] n77;
wire      [7:0] n78;
wire      [7:0] n79;
wire      [7:0] n80;
wire      [7:0] n81;
wire      [7:0] n82;
wire      [7:0] n83;
wire      [7:0] n84;
wire     [15:0] n85;
wire     [23:0] n86;
wire     [31:0] n87;
wire     [39:0] n88;
wire     [47:0] n89;
wire     [55:0] n90;
wire     [63:0] n91;
wire     [71:0] n92;
wire      [7:0] n93;
wire      [7:0] n94;
wire      [7:0] n95;
wire      [7:0] n96;
wire      [7:0] n97;
wire      [7:0] n98;
wire      [7:0] n99;
wire      [7:0] n100;
wire      [7:0] n101;
wire     [15:0] n102;
wire     [23:0] n103;
wire     [31:0] n104;
wire     [39:0] n105;
wire     [47:0] n106;
wire     [55:0] n107;
wire     [63:0] n108;
wire     [71:0] n109;
wire      [7:0] n110;
wire      [7:0] n111;
wire      [7:0] n112;
wire      [7:0] n113;
wire      [7:0] n114;
wire      [7:0] n115;
wire      [7:0] n116;
wire      [7:0] n117;
wire      [7:0] n118;
wire     [15:0] n119;
wire     [23:0] n120;
wire     [31:0] n121;
wire     [39:0] n122;
wire     [47:0] n123;
wire     [55:0] n124;
wire     [63:0] n125;
wire     [71:0] n126;
wire      [7:0] n127;
wire      [7:0] n128;
wire      [7:0] n129;
wire      [7:0] n130;
wire      [7:0] n131;
wire      [7:0] n132;
wire      [7:0] n133;
wire      [7:0] n134;
wire      [7:0] n135;
wire     [15:0] n136;
wire     [23:0] n137;
wire     [31:0] n138;
wire     [39:0] n139;
wire     [47:0] n140;
wire     [55:0] n141;
wire     [63:0] n142;
wire     [71:0] n143;
wire      [7:0] n144;
wire      [7:0] n145;
wire      [7:0] n146;
wire      [7:0] n147;
wire      [7:0] n148;
wire      [7:0] n149;
wire      [7:0] n150;
wire      [7:0] n151;
wire      [7:0] n152;
wire     [15:0] n153;
wire     [23:0] n154;
wire     [31:0] n155;
wire     [39:0] n156;
wire     [47:0] n157;
wire     [55:0] n158;
wire     [63:0] n159;
wire     [71:0] n160;
wire      [7:0] n161;
wire      [7:0] n162;
wire      [7:0] n163;
wire      [7:0] n164;
wire      [7:0] n165;
wire      [7:0] n166;
wire      [7:0] n167;
wire      [7:0] n168;
wire      [7:0] n169;
wire     [15:0] n170;
wire     [23:0] n171;
wire     [31:0] n172;
wire     [39:0] n173;
wire     [47:0] n174;
wire     [55:0] n175;
wire     [63:0] n176;
wire     [71:0] n177;
wire      [7:0] n178;
wire      [7:0] n179;
wire      [7:0] n180;
wire      [7:0] n181;
wire      [7:0] n182;
wire      [7:0] n183;
wire      [7:0] n184;
wire      [7:0] n185;
wire      [7:0] n186;
wire     [15:0] n187;
wire     [23:0] n188;
wire     [31:0] n189;
wire     [39:0] n190;
wire     [47:0] n191;
wire     [55:0] n192;
wire     [63:0] n193;
wire     [71:0] n194;
wire      [7:0] n195;
wire      [7:0] n196;
wire      [7:0] n197;
wire      [7:0] n198;
wire      [7:0] n199;
wire      [7:0] n200;
wire      [7:0] n201;
wire      [7:0] n202;
wire      [7:0] n203;
wire     [15:0] n204;
wire     [23:0] n205;
wire     [31:0] n206;
wire     [39:0] n207;
wire     [47:0] n208;
wire     [55:0] n209;
wire     [63:0] n210;
wire     [71:0] n211;
wire    [143:0] n212;
wire    [215:0] n213;
wire    [287:0] n214;
wire    [359:0] n215;
wire    [431:0] n216;
wire    [503:0] n217;
wire    [575:0] n218;
wire    [647:0] n219;
wire    [647:0] n220;
wire    [647:0] n221;
wire      [7:0] n222;
wire      [7:0] n223;
wire      [7:0] n224;
wire      [7:0] n225;
wire      [7:0] n226;
wire      [7:0] n227;
wire      [7:0] n228;
wire            n229;
wire            n230;
wire            n231;
wire            n232;
wire            n233;
wire            n234;
wire            n235;
wire            n236;
wire            n237;
wire            n238;
wire            n239;
wire      [8:0] n240;
wire            n241;
wire      [9:0] n242;
wire            n243;
wire            n244;
wire            n245;
wire            n246;
wire            n247;
wire            n248;
wire            n249;
wire            n250;
wire            n251;
wire            n252;
wire      [7:0] n253;
wire      [7:0] n254;
wire      [7:0] n255;
wire      [7:0] n256;
wire      [7:0] n257;
wire            n258;
wire      [3:0] n259;
wire      [3:0] n260;
wire      [3:0] n261;
wire      [7:0] n262;
wire      [7:0] n263;
wire      [7:0] n264;
wire    [647:0] n265;
wire    [647:0] n266;
wire    [647:0] n267;
wire            n268;
wire            n269;
wire            n270;
wire     [71:0] n271;
wire     [71:0] n272;
wire     [71:0] n273;
wire     [71:0] n274;
wire     [71:0] n275;
wire     [71:0] n276;
wire     [71:0] n277;
wire     [71:0] n278;
wire     [71:0] n279;
wire     [71:0] n280;
wire     [71:0] n281;
wire     [71:0] n282;
wire     [71:0] n283;
wire     [71:0] n284;
wire     [71:0] n285;
wire     [71:0] n286;
wire     [71:0] n287;
wire     [71:0] n288;
wire     [71:0] n289;
wire     [71:0] n290;
wire     [71:0] n291;
wire     [71:0] n292;
wire     [71:0] n293;
wire     [71:0] n294;
wire     [71:0] n295;
wire     [71:0] n296;
wire     [71:0] n297;
wire     [71:0] n298;
wire     [71:0] n299;
wire     [71:0] n300;
wire     [71:0] n301;
wire     [71:0] n302;
wire     [71:0] n303;
wire     [71:0] n304;
wire     [71:0] n305;
wire     [71:0] n306;
wire     [71:0] n307;
wire     [71:0] n308;
wire     [71:0] n309;
wire     [71:0] n310;
wire     [71:0] n311;
wire     [71:0] n312;
wire     [71:0] n313;
wire     [71:0] n314;
wire     [71:0] n315;
wire     [71:0] n316;
wire     [71:0] n317;
wire     [71:0] n318;
wire            n319;
wire      [8:0] n320;
wire      [7:0] n321;
wire            n322;
wire      [7:0] n323;
wire            n324;
wire      [7:0] n325;
wire            n326;
wire      [7:0] n327;
wire            n328;
wire      [7:0] n329;
wire            n330;
wire      [7:0] n331;
wire            n332;
wire      [7:0] n333;
wire      [7:0] n334;
wire      [7:0] n335;
wire      [7:0] n336;
wire      [7:0] n337;
wire      [7:0] n338;
wire      [7:0] n339;
wire      [7:0] n340;
wire      [7:0] n341;
wire      [7:0] n342;
wire      [7:0] n343;
wire      [7:0] n344;
wire      [7:0] n345;
wire      [7:0] n346;
wire      [7:0] n347;
wire      [7:0] n348;
wire      [7:0] n349;
wire      [7:0] n350;
wire      [7:0] n351;
wire      [7:0] n352;
wire      [7:0] n353;
wire      [7:0] n354;
wire      [7:0] n355;
wire      [7:0] n356;
wire      [7:0] n357;
wire      [7:0] n358;
wire      [7:0] n359;
wire      [7:0] n360;
wire      [7:0] n361;
wire      [7:0] n362;
wire      [7:0] n363;
wire      [7:0] n364;
wire      [7:0] n365;
wire      [7:0] n366;
wire      [7:0] n367;
wire      [7:0] n368;
wire      [7:0] n369;
wire      [7:0] n370;
wire      [7:0] n371;
wire      [7:0] n372;
wire      [7:0] n373;
wire      [7:0] n374;
wire      [7:0] n375;
wire      [7:0] n376;
wire      [7:0] n377;
wire      [7:0] n378;
wire      [7:0] n379;
wire      [7:0] n380;
wire      [7:0] n381;
wire      [7:0] n382;
wire      [7:0] n383;
wire      [7:0] n384;
wire      [7:0] n385;
wire      [7:0] n386;
wire      [7:0] n387;
wire      [7:0] n388;
wire      [7:0] n389;
wire      [7:0] n390;
wire     [15:0] n391;
wire     [23:0] n392;
wire     [31:0] n393;
wire     [39:0] n394;
wire     [47:0] n395;
wire     [55:0] n396;
wire     [63:0] n397;
wire     [71:0] n398;
wire     [71:0] n399;
wire     [71:0] n400;
wire     [71:0] n401;
wire     [71:0] n402;
wire     [71:0] n403;
wire     [71:0] n404;
wire      [8:0] RAM_0_addr0;
wire      [7:0] RAM_0_data0;
wire            n405;
wire            n406;
wire            n407;
wire            n408;
wire            n409;
wire            n410;
wire            n411;
wire            n412;
wire            n413;
wire            n414;
wire            n415;
wire            n416;
wire            n417;
wire            n418;
wire            n419;
wire            n420;
wire      [8:0] RAM_1_addr0;
wire      [7:0] RAM_1_data0;
wire            n421;
wire            n422;
wire            n423;
wire      [8:0] RAM_2_addr0;
wire      [7:0] RAM_2_data0;
wire            n424;
wire            n425;
wire            n426;
wire      [8:0] RAM_3_addr0;
wire      [7:0] RAM_3_data0;
wire            n427;
wire            n428;
wire            n429;
wire      [8:0] RAM_4_addr0;
wire      [7:0] RAM_4_data0;
wire            n430;
wire            n431;
wire            n432;
wire      [8:0] RAM_5_addr0;
wire      [7:0] RAM_5_data0;
wire            n433;
wire            n434;
wire            n435;
wire      [8:0] RAM_6_addr0;
wire      [7:0] RAM_6_data0;
wire            n436;
wire            n437;
wire            n438;
wire      [8:0] RAM_7_addr0;
wire      [7:0] RAM_7_data0;
wire            n439;
wire            n440;
wire            n441;
reg      [7:0] RAM_0[511:0];
reg      [7:0] RAM_1[511:0];
reg      [7:0] RAM_2[511:0];
reg      [7:0] RAM_3[511:0];
reg      [7:0] RAM_4[511:0];
reg      [7:0] RAM_5[511:0];
reg      [7:0] RAM_6[511:0];
reg      [7:0] RAM_7[511:0];
wire clk;
wire rst;
wire step;
assign n0 =  ( arg_1_TVALID ) == ( 1'd0 )  ;
assign n1 =  ( arg_0_TVALID ) == ( 1'd1 )  ;
assign n2 =  ( n0 ) & ( n1 )  ;
assign n3 =  ( arg_0_TREADY ) == ( 1'd1 )  ;
assign n4 =  ( n2 ) & ( n3 )  ;
assign n5 =  ( arg_1_TREADY ) == ( 1'd0 )  ;
assign n6 =  ( arg_0_TREADY ) == ( 1'd0 )  ;
assign n7 =  ( n5 ) & ( n6 )  ;
assign n8 =  ( st_ready ) == ( 1'd0 )  ;
assign n9 =  ( n7 ) & ( n8 )  ;
assign n10 =  ( st_ready ) == ( 1'd1 )  ;
assign n11 =  ( n7 ) & ( n10 )  ;
assign n12 =  ( RAM_x ) == ( 9'd0 )  ;
assign n13 =  ( n11 ) & ( n12 )  ;
assign n14 =  ( RAM_y ) == ( 10'd0 )  ;
assign n15 =  ( n13 ) & ( n14 )  ;
assign n16 =  ( n12 ) & ( n14 )  ;
assign n17 = ~ ( n16 ) ;
assign n18 =  ( n11 ) & ( n17 )  ;
assign n19 =  ( RAM_x ) == ( 9'd488 )  ;
assign n20 =  ( RAM_w ) == ( 3'd7 )  ;
assign n21 =  ( RAM_w ) + ( 3'd1 )  ;
assign n22 =  ( n20 ) ? ( 3'd0 ) : ( n21 ) ;
assign n23 =  ( n19 ) ? ( n22 ) : ( RAM_w ) ;
assign n24 =  ( arg_1_TVALID ) == ( 1'd1 )  ;
assign n25 =  ( arg_1_TREADY ) == ( 1'd1 )  ;
assign n26 =  ( n24 ) & ( n25 )  ;
assign n27 =  ( arg_0_TVALID ) == ( 1'd0 )  ;
assign n28 =  ( n26 ) & ( n27 )  ;
assign n29 =  ( n28 ) & ( n6 )  ;
assign n30 =  ( n29 ) ? ( RAM_w ) : ( RAM_w ) ;
assign n31 =  ( n18 ) ? ( n23 ) : ( n30 ) ;
assign n32 =  ( n15 ) ? ( RAM_w ) : ( n31 ) ;
assign n33 =  ( n9 ) ? ( RAM_w ) : ( n32 ) ;
assign n34 =  ( n4 ) ? ( RAM_w ) : ( n33 ) ;
assign n35 =  ( RAM_x ) + ( 9'd1 )  ;
assign n36 =  ( n19 ) ? ( 9'd1 ) : ( n35 ) ;
assign n37 =  ( n29 ) ? ( RAM_x ) : ( RAM_x ) ;
assign n38 =  ( n18 ) ? ( n36 ) : ( n37 ) ;
assign n39 =  ( n15 ) ? ( 9'd1 ) : ( n38 ) ;
assign n40 =  ( n9 ) ? ( RAM_x ) : ( n39 ) ;
assign n41 =  ( n4 ) ? ( RAM_x ) : ( n40 ) ;
assign n42 =  ( RAM_y ) == ( 10'd648 )  ;
assign n43 =  ( RAM_y ) + ( 10'd1 )  ;
assign n44 =  ( n42 ) ? ( 10'd0 ) : ( n43 ) ;
assign n45 =  ( n19 ) ? ( n44 ) : ( RAM_y ) ;
assign n46 =  ( n29 ) ? ( RAM_y ) : ( RAM_y ) ;
assign n47 =  ( n18 ) ? ( n45 ) : ( n46 ) ;
assign n48 =  ( n15 ) ? ( RAM_y ) : ( n47 ) ;
assign n49 =  ( n9 ) ? ( RAM_y ) : ( n48 ) ;
assign n50 =  ( n4 ) ? ( RAM_y ) : ( n49 ) ;
assign n51 =  ( RAM_x ) == ( 9'd1 )  ;
assign n52 =  ( n51 ) & ( n42 )  ;
assign n53 =  ( RAM_x ) > ( 9'd8 )  ;
assign n54 =  ( RAM_y ) >= ( 10'd8 )  ;
assign n55 =  ( n53 ) & ( n54 )  ;
assign n56 =  ( RAM_y ) > ( 10'd8 )  ;
assign n57 =  ( n51 ) & ( n56 )  ;
assign n58 =  ( n55 ) | ( n57 )  ;
assign n59 = stencil_8[71:64] ;
assign n60 = stencil_7[71:64] ;
assign n61 = stencil_6[71:64] ;
assign n62 = stencil_5[71:64] ;
assign n63 = stencil_4[71:64] ;
assign n64 = stencil_3[71:64] ;
assign n65 = stencil_2[71:64] ;
assign n66 = stencil_1[71:64] ;
assign n67 = stencil_0[71:64] ;
assign n68 =  { ( n66 ) , ( n67 ) }  ;
assign n69 =  { ( n65 ) , ( n68 ) }  ;
assign n70 =  { ( n64 ) , ( n69 ) }  ;
assign n71 =  { ( n63 ) , ( n70 ) }  ;
assign n72 =  { ( n62 ) , ( n71 ) }  ;
assign n73 =  { ( n61 ) , ( n72 ) }  ;
assign n74 =  { ( n60 ) , ( n73 ) }  ;
assign n75 =  { ( n59 ) , ( n74 ) }  ;
assign n76 = stencil_8[63:56] ;
assign n77 = stencil_7[63:56] ;
assign n78 = stencil_6[63:56] ;
assign n79 = stencil_5[63:56] ;
assign n80 = stencil_4[63:56] ;
assign n81 = stencil_3[63:56] ;
assign n82 = stencil_2[63:56] ;
assign n83 = stencil_1[63:56] ;
assign n84 = stencil_0[63:56] ;
assign n85 =  { ( n83 ) , ( n84 ) }  ;
assign n86 =  { ( n82 ) , ( n85 ) }  ;
assign n87 =  { ( n81 ) , ( n86 ) }  ;
assign n88 =  { ( n80 ) , ( n87 ) }  ;
assign n89 =  { ( n79 ) , ( n88 ) }  ;
assign n90 =  { ( n78 ) , ( n89 ) }  ;
assign n91 =  { ( n77 ) , ( n90 ) }  ;
assign n92 =  { ( n76 ) , ( n91 ) }  ;
assign n93 = stencil_8[55:48] ;
assign n94 = stencil_7[55:48] ;
assign n95 = stencil_6[55:48] ;
assign n96 = stencil_5[55:48] ;
assign n97 = stencil_4[55:48] ;
assign n98 = stencil_3[55:48] ;
assign n99 = stencil_2[55:48] ;
assign n100 = stencil_1[55:48] ;
assign n101 = stencil_0[55:48] ;
assign n102 =  { ( n100 ) , ( n101 ) }  ;
assign n103 =  { ( n99 ) , ( n102 ) }  ;
assign n104 =  { ( n98 ) , ( n103 ) }  ;
assign n105 =  { ( n97 ) , ( n104 ) }  ;
assign n106 =  { ( n96 ) , ( n105 ) }  ;
assign n107 =  { ( n95 ) , ( n106 ) }  ;
assign n108 =  { ( n94 ) , ( n107 ) }  ;
assign n109 =  { ( n93 ) , ( n108 ) }  ;
assign n110 = stencil_8[47:40] ;
assign n111 = stencil_7[47:40] ;
assign n112 = stencil_6[47:40] ;
assign n113 = stencil_5[47:40] ;
assign n114 = stencil_4[47:40] ;
assign n115 = stencil_3[47:40] ;
assign n116 = stencil_2[47:40] ;
assign n117 = stencil_1[47:40] ;
assign n118 = stencil_0[47:40] ;
assign n119 =  { ( n117 ) , ( n118 ) }  ;
assign n120 =  { ( n116 ) , ( n119 ) }  ;
assign n121 =  { ( n115 ) , ( n120 ) }  ;
assign n122 =  { ( n114 ) , ( n121 ) }  ;
assign n123 =  { ( n113 ) , ( n122 ) }  ;
assign n124 =  { ( n112 ) , ( n123 ) }  ;
assign n125 =  { ( n111 ) , ( n124 ) }  ;
assign n126 =  { ( n110 ) , ( n125 ) }  ;
assign n127 = stencil_8[39:32] ;
assign n128 = stencil_7[39:32] ;
assign n129 = stencil_6[39:32] ;
assign n130 = stencil_5[39:32] ;
assign n131 = stencil_4[39:32] ;
assign n132 = stencil_3[39:32] ;
assign n133 = stencil_2[39:32] ;
assign n134 = stencil_1[39:32] ;
assign n135 = stencil_0[39:32] ;
assign n136 =  { ( n134 ) , ( n135 ) }  ;
assign n137 =  { ( n133 ) , ( n136 ) }  ;
assign n138 =  { ( n132 ) , ( n137 ) }  ;
assign n139 =  { ( n131 ) , ( n138 ) }  ;
assign n140 =  { ( n130 ) , ( n139 ) }  ;
assign n141 =  { ( n129 ) , ( n140 ) }  ;
assign n142 =  { ( n128 ) , ( n141 ) }  ;
assign n143 =  { ( n127 ) , ( n142 ) }  ;
assign n144 = stencil_8[31:24] ;
assign n145 = stencil_7[31:24] ;
assign n146 = stencil_6[31:24] ;
assign n147 = stencil_5[31:24] ;
assign n148 = stencil_4[31:24] ;
assign n149 = stencil_3[31:24] ;
assign n150 = stencil_2[31:24] ;
assign n151 = stencil_1[31:24] ;
assign n152 = stencil_0[31:24] ;
assign n153 =  { ( n151 ) , ( n152 ) }  ;
assign n154 =  { ( n150 ) , ( n153 ) }  ;
assign n155 =  { ( n149 ) , ( n154 ) }  ;
assign n156 =  { ( n148 ) , ( n155 ) }  ;
assign n157 =  { ( n147 ) , ( n156 ) }  ;
assign n158 =  { ( n146 ) , ( n157 ) }  ;
assign n159 =  { ( n145 ) , ( n158 ) }  ;
assign n160 =  { ( n144 ) , ( n159 ) }  ;
assign n161 = stencil_8[23:16] ;
assign n162 = stencil_7[23:16] ;
assign n163 = stencil_6[23:16] ;
assign n164 = stencil_5[23:16] ;
assign n165 = stencil_4[23:16] ;
assign n166 = stencil_3[23:16] ;
assign n167 = stencil_2[23:16] ;
assign n168 = stencil_1[23:16] ;
assign n169 = stencil_0[23:16] ;
assign n170 =  { ( n168 ) , ( n169 ) }  ;
assign n171 =  { ( n167 ) , ( n170 ) }  ;
assign n172 =  { ( n166 ) , ( n171 ) }  ;
assign n173 =  { ( n165 ) , ( n172 ) }  ;
assign n174 =  { ( n164 ) , ( n173 ) }  ;
assign n175 =  { ( n163 ) , ( n174 ) }  ;
assign n176 =  { ( n162 ) , ( n175 ) }  ;
assign n177 =  { ( n161 ) , ( n176 ) }  ;
assign n178 = stencil_8[15:8] ;
assign n179 = stencil_7[15:8] ;
assign n180 = stencil_6[15:8] ;
assign n181 = stencil_5[15:8] ;
assign n182 = stencil_4[15:8] ;
assign n183 = stencil_3[15:8] ;
assign n184 = stencil_2[15:8] ;
assign n185 = stencil_1[15:8] ;
assign n186 = stencil_0[15:8] ;
assign n187 =  { ( n185 ) , ( n186 ) }  ;
assign n188 =  { ( n184 ) , ( n187 ) }  ;
assign n189 =  { ( n183 ) , ( n188 ) }  ;
assign n190 =  { ( n182 ) , ( n189 ) }  ;
assign n191 =  { ( n181 ) , ( n190 ) }  ;
assign n192 =  { ( n180 ) , ( n191 ) }  ;
assign n193 =  { ( n179 ) , ( n192 ) }  ;
assign n194 =  { ( n178 ) , ( n193 ) }  ;
assign n195 = stencil_8[7:0] ;
assign n196 = stencil_7[7:0] ;
assign n197 = stencil_6[7:0] ;
assign n198 = stencil_5[7:0] ;
assign n199 = stencil_4[7:0] ;
assign n200 = stencil_3[7:0] ;
assign n201 = stencil_2[7:0] ;
assign n202 = stencil_1[7:0] ;
assign n203 = stencil_0[7:0] ;
assign n204 =  { ( n202 ) , ( n203 ) }  ;
assign n205 =  { ( n201 ) , ( n204 ) }  ;
assign n206 =  { ( n200 ) , ( n205 ) }  ;
assign n207 =  { ( n199 ) , ( n206 ) }  ;
assign n208 =  { ( n198 ) , ( n207 ) }  ;
assign n209 =  { ( n197 ) , ( n208 ) }  ;
assign n210 =  { ( n196 ) , ( n209 ) }  ;
assign n211 =  { ( n195 ) , ( n210 ) }  ;
assign n212 =  { ( n194 ) , ( n211 ) }  ;
assign n213 =  { ( n177 ) , ( n212 ) }  ;
assign n214 =  { ( n160 ) , ( n213 ) }  ;
assign n215 =  { ( n143 ) , ( n214 ) }  ;
assign n216 =  { ( n126 ) , ( n215 ) }  ;
assign n217 =  { ( n109 ) , ( n216 ) }  ;
assign n218 =  { ( n92 ) , ( n217 ) }  ;
assign n219 =  { ( n75 ) , ( n218 ) }  ;
assign n220 =  ( n58 ) ? ( n219 ) : ( proc_in ) ;
assign n221 =  ( n52 ) ? ( proc_in ) : ( n220 ) ;
assign n222 = gb_fun(n221) ;
assign n223 =  ( n52 ) ? ( arg_0_TDATA ) : ( n222 ) ;
assign n224 =  ( n29 ) ? ( arg_0_TDATA ) : ( arg_0_TDATA ) ;
assign n225 =  ( n18 ) ? ( arg_0_TDATA ) : ( n224 ) ;
assign n226 =  ( n15 ) ? ( arg_0_TDATA ) : ( n225 ) ;
assign n227 =  ( n9 ) ? ( n223 ) : ( n226 ) ;
assign n228 =  ( n4 ) ? ( arg_0_TDATA ) : ( n227 ) ;
assign n229 =  ( gbit ) == ( 4'd0 )  ;
assign n230 =  ( gbit ) == ( 4'd7 )  ;
assign n231 =  ( n229 ) | ( n230 )  ;
assign n232 =  ( n231 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n233 =  ( n58 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n234 =  ( n52 ) ? ( arg_0_TVALID ) : ( n233 ) ;
assign n235 =  ( n29 ) ? ( 1'd0 ) : ( arg_0_TVALID ) ;
assign n236 =  ( n18 ) ? ( arg_0_TVALID ) : ( n235 ) ;
assign n237 =  ( n15 ) ? ( 1'd0 ) : ( n236 ) ;
assign n238 =  ( n9 ) ? ( n234 ) : ( n237 ) ;
assign n239 =  ( n4 ) ? ( n232 ) : ( n238 ) ;
assign n240 =  ( 9'd488 ) - ( 9'd1 )  ;
assign n241 =  ( RAM_x ) == ( n240 )  ;
assign n242 =  ( 10'd648 ) - ( 10'd1 )  ;
assign n243 =  ( RAM_y ) == ( n242 )  ;
assign n244 =  ( n241 ) & ( n243 )  ;
assign n245 =  ( n244 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n246 =  ( RAM_y ) < ( 10'd8 )  ;
assign n247 =  ( n246 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n248 =  ( n29 ) ? ( 1'd0 ) : ( arg_1_TREADY ) ;
assign n249 =  ( n18 ) ? ( n247 ) : ( n248 ) ;
assign n250 =  ( n15 ) ? ( 1'd1 ) : ( n249 ) ;
assign n251 =  ( n9 ) ? ( n245 ) : ( n250 ) ;
assign n252 =  ( n4 ) ? ( arg_1_TREADY ) : ( n251 ) ;
assign n253 =  ( n29 ) ? ( arg_1_TDATA ) : ( cur_pix ) ;
assign n254 =  ( n18 ) ? ( cur_pix ) : ( n253 ) ;
assign n255 =  ( n15 ) ? ( cur_pix ) : ( n254 ) ;
assign n256 =  ( n9 ) ? ( cur_pix ) : ( n255 ) ;
assign n257 =  ( n4 ) ? ( cur_pix ) : ( n256 ) ;
assign n258 =  ( n19 ) & ( n42 )  ;
assign n259 =  ( gbit ) + ( 4'd1 )  ;
assign n260 =  ( n258 ) ? ( n259 ) : ( gbit ) ;
assign n261 =  ( n4 ) ? ( n260 ) : ( gbit ) ;
assign n262 =  ( n18 ) ? ( cur_pix ) : ( pre_pix ) ;
assign n263 =  ( n15 ) ? ( cur_pix ) : ( n262 ) ;
assign n264 =  ( n9 ) ? ( pre_pix ) : ( n263 ) ;
assign n265 =  ( n18 ) ? ( proc_in ) : ( proc_in ) ;
assign n266 =  ( n15 ) ? ( proc_in ) : ( n265 ) ;
assign n267 =  ( n9 ) ? ( n221 ) : ( n266 ) ;
assign n268 =  ( n18 ) ? ( n247 ) : ( st_ready ) ;
assign n269 =  ( n15 ) ? ( 1'd1 ) : ( n268 ) ;
assign n270 =  ( n9 ) ? ( 1'd1 ) : ( n269 ) ;
assign n271 =  ( n246 ) ? ( stencil_0 ) : ( stencil_1 ) ;
assign n272 =  ( n29 ) ? ( stencil_0 ) : ( stencil_0 ) ;
assign n273 =  ( n18 ) ? ( stencil_0 ) : ( n272 ) ;
assign n274 =  ( n15 ) ? ( stencil_0 ) : ( n273 ) ;
assign n275 =  ( n9 ) ? ( n271 ) : ( n274 ) ;
assign n276 =  ( n4 ) ? ( stencil_0 ) : ( n275 ) ;
assign n277 =  ( n246 ) ? ( stencil_1 ) : ( stencil_2 ) ;
assign n278 =  ( n29 ) ? ( stencil_1 ) : ( stencil_1 ) ;
assign n279 =  ( n18 ) ? ( stencil_1 ) : ( n278 ) ;
assign n280 =  ( n15 ) ? ( stencil_1 ) : ( n279 ) ;
assign n281 =  ( n9 ) ? ( n277 ) : ( n280 ) ;
assign n282 =  ( n4 ) ? ( stencil_1 ) : ( n281 ) ;
assign n283 =  ( n246 ) ? ( stencil_2 ) : ( stencil_3 ) ;
assign n284 =  ( n29 ) ? ( stencil_2 ) : ( stencil_2 ) ;
assign n285 =  ( n18 ) ? ( stencil_2 ) : ( n284 ) ;
assign n286 =  ( n15 ) ? ( stencil_2 ) : ( n285 ) ;
assign n287 =  ( n9 ) ? ( n283 ) : ( n286 ) ;
assign n288 =  ( n4 ) ? ( stencil_2 ) : ( n287 ) ;
assign n289 =  ( n246 ) ? ( stencil_3 ) : ( stencil_4 ) ;
assign n290 =  ( n29 ) ? ( stencil_3 ) : ( stencil_3 ) ;
assign n291 =  ( n18 ) ? ( stencil_3 ) : ( n290 ) ;
assign n292 =  ( n15 ) ? ( stencil_3 ) : ( n291 ) ;
assign n293 =  ( n9 ) ? ( n289 ) : ( n292 ) ;
assign n294 =  ( n4 ) ? ( stencil_3 ) : ( n293 ) ;
assign n295 =  ( n246 ) ? ( stencil_4 ) : ( stencil_5 ) ;
assign n296 =  ( n29 ) ? ( stencil_4 ) : ( stencil_4 ) ;
assign n297 =  ( n18 ) ? ( stencil_4 ) : ( n296 ) ;
assign n298 =  ( n15 ) ? ( stencil_4 ) : ( n297 ) ;
assign n299 =  ( n9 ) ? ( n295 ) : ( n298 ) ;
assign n300 =  ( n4 ) ? ( stencil_4 ) : ( n299 ) ;
assign n301 =  ( n246 ) ? ( stencil_5 ) : ( stencil_6 ) ;
assign n302 =  ( n29 ) ? ( stencil_5 ) : ( stencil_5 ) ;
assign n303 =  ( n18 ) ? ( stencil_5 ) : ( n302 ) ;
assign n304 =  ( n15 ) ? ( stencil_5 ) : ( n303 ) ;
assign n305 =  ( n9 ) ? ( n301 ) : ( n304 ) ;
assign n306 =  ( n4 ) ? ( stencil_5 ) : ( n305 ) ;
assign n307 =  ( n246 ) ? ( stencil_6 ) : ( stencil_7 ) ;
assign n308 =  ( n29 ) ? ( stencil_6 ) : ( stencil_6 ) ;
assign n309 =  ( n18 ) ? ( stencil_6 ) : ( n308 ) ;
assign n310 =  ( n15 ) ? ( stencil_6 ) : ( n309 ) ;
assign n311 =  ( n9 ) ? ( n307 ) : ( n310 ) ;
assign n312 =  ( n4 ) ? ( stencil_6 ) : ( n311 ) ;
assign n313 =  ( n246 ) ? ( stencil_7 ) : ( stencil_8 ) ;
assign n314 =  ( n29 ) ? ( stencil_7 ) : ( stencil_7 ) ;
assign n315 =  ( n18 ) ? ( stencil_7 ) : ( n314 ) ;
assign n316 =  ( n15 ) ? ( stencil_7 ) : ( n315 ) ;
assign n317 =  ( n9 ) ? ( n313 ) : ( n316 ) ;
assign n318 =  ( n4 ) ? ( stencil_7 ) : ( n317 ) ;
assign n319 =  ( RAM_w ) == ( 3'd0 )  ;
assign n320 =  ( RAM_x ) - ( 9'd1 )  ;
assign n321 =  (  RAM_7 [ n320 ] )  ;
assign n322 =  ( RAM_w ) == ( 3'd1 )  ;
assign n323 =  (  RAM_0 [ n320 ] )  ;
assign n324 =  ( RAM_w ) == ( 3'd2 )  ;
assign n325 =  (  RAM_1 [ n320 ] )  ;
assign n326 =  ( RAM_w ) == ( 3'd3 )  ;
assign n327 =  (  RAM_2 [ n320 ] )  ;
assign n328 =  ( RAM_w ) == ( 3'd4 )  ;
assign n329 =  (  RAM_3 [ n320 ] )  ;
assign n330 =  ( RAM_w ) == ( 3'd5 )  ;
assign n331 =  (  RAM_4 [ n320 ] )  ;
assign n332 =  ( RAM_w ) == ( 3'd6 )  ;
assign n333 =  (  RAM_5 [ n320 ] )  ;
assign n334 =  (  RAM_6 [ n320 ] )  ;
assign n335 =  ( n332 ) ? ( n333 ) : ( n334 ) ;
assign n336 =  ( n330 ) ? ( n331 ) : ( n335 ) ;
assign n337 =  ( n328 ) ? ( n329 ) : ( n336 ) ;
assign n338 =  ( n326 ) ? ( n327 ) : ( n337 ) ;
assign n339 =  ( n324 ) ? ( n325 ) : ( n338 ) ;
assign n340 =  ( n322 ) ? ( n323 ) : ( n339 ) ;
assign n341 =  ( n319 ) ? ( n321 ) : ( n340 ) ;
assign n342 =  ( n332 ) ? ( n331 ) : ( n333 ) ;
assign n343 =  ( n330 ) ? ( n329 ) : ( n342 ) ;
assign n344 =  ( n328 ) ? ( n327 ) : ( n343 ) ;
assign n345 =  ( n326 ) ? ( n325 ) : ( n344 ) ;
assign n346 =  ( n324 ) ? ( n323 ) : ( n345 ) ;
assign n347 =  ( n322 ) ? ( n321 ) : ( n346 ) ;
assign n348 =  ( n319 ) ? ( n334 ) : ( n347 ) ;
assign n349 =  ( n332 ) ? ( n329 ) : ( n331 ) ;
assign n350 =  ( n330 ) ? ( n327 ) : ( n349 ) ;
assign n351 =  ( n328 ) ? ( n325 ) : ( n350 ) ;
assign n352 =  ( n326 ) ? ( n323 ) : ( n351 ) ;
assign n353 =  ( n324 ) ? ( n321 ) : ( n352 ) ;
assign n354 =  ( n322 ) ? ( n334 ) : ( n353 ) ;
assign n355 =  ( n319 ) ? ( n333 ) : ( n354 ) ;
assign n356 =  ( n332 ) ? ( n327 ) : ( n329 ) ;
assign n357 =  ( n330 ) ? ( n325 ) : ( n356 ) ;
assign n358 =  ( n328 ) ? ( n323 ) : ( n357 ) ;
assign n359 =  ( n326 ) ? ( n321 ) : ( n358 ) ;
assign n360 =  ( n324 ) ? ( n334 ) : ( n359 ) ;
assign n361 =  ( n322 ) ? ( n333 ) : ( n360 ) ;
assign n362 =  ( n319 ) ? ( n331 ) : ( n361 ) ;
assign n363 =  ( n332 ) ? ( n325 ) : ( n327 ) ;
assign n364 =  ( n330 ) ? ( n323 ) : ( n363 ) ;
assign n365 =  ( n328 ) ? ( n321 ) : ( n364 ) ;
assign n366 =  ( n326 ) ? ( n334 ) : ( n365 ) ;
assign n367 =  ( n324 ) ? ( n333 ) : ( n366 ) ;
assign n368 =  ( n322 ) ? ( n331 ) : ( n367 ) ;
assign n369 =  ( n319 ) ? ( n329 ) : ( n368 ) ;
assign n370 =  ( n332 ) ? ( n323 ) : ( n325 ) ;
assign n371 =  ( n330 ) ? ( n321 ) : ( n370 ) ;
assign n372 =  ( n328 ) ? ( n334 ) : ( n371 ) ;
assign n373 =  ( n326 ) ? ( n333 ) : ( n372 ) ;
assign n374 =  ( n324 ) ? ( n331 ) : ( n373 ) ;
assign n375 =  ( n322 ) ? ( n329 ) : ( n374 ) ;
assign n376 =  ( n319 ) ? ( n327 ) : ( n375 ) ;
assign n377 =  ( n332 ) ? ( n321 ) : ( n323 ) ;
assign n378 =  ( n330 ) ? ( n334 ) : ( n377 ) ;
assign n379 =  ( n328 ) ? ( n333 ) : ( n378 ) ;
assign n380 =  ( n326 ) ? ( n331 ) : ( n379 ) ;
assign n381 =  ( n324 ) ? ( n329 ) : ( n380 ) ;
assign n382 =  ( n322 ) ? ( n327 ) : ( n381 ) ;
assign n383 =  ( n319 ) ? ( n325 ) : ( n382 ) ;
assign n384 =  ( n332 ) ? ( n334 ) : ( n321 ) ;
assign n385 =  ( n330 ) ? ( n333 ) : ( n384 ) ;
assign n386 =  ( n328 ) ? ( n331 ) : ( n385 ) ;
assign n387 =  ( n326 ) ? ( n329 ) : ( n386 ) ;
assign n388 =  ( n324 ) ? ( n327 ) : ( n387 ) ;
assign n389 =  ( n322 ) ? ( n325 ) : ( n388 ) ;
assign n390 =  ( n319 ) ? ( n323 ) : ( n389 ) ;
assign n391 =  { ( n383 ) , ( n390 ) }  ;
assign n392 =  { ( n376 ) , ( n391 ) }  ;
assign n393 =  { ( n369 ) , ( n392 ) }  ;
assign n394 =  { ( n362 ) , ( n393 ) }  ;
assign n395 =  { ( n355 ) , ( n394 ) }  ;
assign n396 =  { ( n348 ) , ( n395 ) }  ;
assign n397 =  { ( n341 ) , ( n396 ) }  ;
assign n398 =  { ( pre_pix ) , ( n397 ) }  ;
assign n399 =  ( n246 ) ? ( stencil_8 ) : ( n398 ) ;
assign n400 =  ( n29 ) ? ( stencil_8 ) : ( stencil_8 ) ;
assign n401 =  ( n18 ) ? ( n399 ) : ( n400 ) ;
assign n402 =  ( n15 ) ? ( stencil_8 ) : ( n401 ) ;
assign n403 =  ( n9 ) ? ( stencil_8 ) : ( n402 ) ;
assign n404 =  ( n4 ) ? ( stencil_8 ) : ( n403 ) ;
assign n405 = ~ ( n4 ) ;
assign n406 = ~ ( n9 ) ;
assign n407 =  ( n405 ) & ( n406 )  ;
assign n408 = ~ ( n15 ) ;
assign n409 =  ( n407 ) & ( n408 )  ;
assign n410 = ~ ( n18 ) ;
assign n411 =  ( n409 ) & ( n410 )  ;
assign n412 = ~ ( n29 ) ;
assign n413 =  ( n411 ) & ( n412 )  ;
assign n414 =  ( n411 ) & ( n29 )  ;
assign n415 =  ( n409 ) & ( n18 )  ;
assign n416 = ~ ( n319 ) ;
assign n417 =  ( n415 ) & ( n416 )  ;
assign n418 =  ( n415 ) & ( n319 )  ;
assign n419 =  ( n407 ) & ( n15 )  ;
assign n420 =  ( n405 ) & ( n9 )  ;
assign RAM_0_addr0 = n418 ? (n320) : (0);
assign RAM_0_data0 = n418 ? (pre_pix) : (RAM_0[0]);
assign n421 = ~ ( n322 ) ;
assign n422 =  ( n415 ) & ( n421 )  ;
assign n423 =  ( n415 ) & ( n322 )  ;
assign RAM_1_addr0 = n423 ? (n320) : (0);
assign RAM_1_data0 = n423 ? (pre_pix) : (RAM_1[0]);
assign n424 = ~ ( n324 ) ;
assign n425 =  ( n415 ) & ( n424 )  ;
assign n426 =  ( n415 ) & ( n324 )  ;
assign RAM_2_addr0 = n426 ? (n320) : (0);
assign RAM_2_data0 = n426 ? (pre_pix) : (RAM_2[0]);
assign n427 = ~ ( n326 ) ;
assign n428 =  ( n415 ) & ( n427 )  ;
assign n429 =  ( n415 ) & ( n326 )  ;
assign RAM_3_addr0 = n429 ? (n320) : (0);
assign RAM_3_data0 = n429 ? (pre_pix) : (RAM_3[0]);
assign n430 = ~ ( n328 ) ;
assign n431 =  ( n415 ) & ( n430 )  ;
assign n432 =  ( n415 ) & ( n328 )  ;
assign RAM_4_addr0 = n432 ? (n320) : (0);
assign RAM_4_data0 = n432 ? (pre_pix) : (RAM_4[0]);
assign n433 = ~ ( n330 ) ;
assign n434 =  ( n415 ) & ( n433 )  ;
assign n435 =  ( n415 ) & ( n330 )  ;
assign RAM_5_addr0 = n435 ? (n320) : (0);
assign RAM_5_data0 = n435 ? (pre_pix) : (RAM_5[0]);
assign n436 = ~ ( n332 ) ;
assign n437 =  ( n415 ) & ( n436 )  ;
assign n438 =  ( n415 ) & ( n332 )  ;
assign RAM_6_addr0 = n438 ? (n320) : (0);
assign RAM_6_data0 = n438 ? (pre_pix) : (RAM_6[0]);
assign n439 = ~ ( n20 ) ;
assign n440 =  ( n415 ) & ( n439 )  ;
assign n441 =  ( n415 ) & ( n20 )  ;
assign RAM_7_addr0 = n441 ? (n320) : (0);
assign RAM_7_data0 = n441 ? (pre_pix) : (RAM_7[0]);
/*
function [7:0] gb_fun ;
input [647:0] arg0;
    begin
//TODO: Add the specific function HERE.    end
endfunction
*/

always @(posedge clk) begin
   if(rst) begin
       RAM_w <= RAM_w;
       RAM_x <= RAM_x;
       RAM_y <= RAM_y;
       arg_0_TDATA <= arg_0_TDATA;
       arg_0_TVALID <= arg_0_TVALID;
       arg_1_TREADY <= arg_1_TREADY;
       cur_pix <= cur_pix;
       gbit <= gbit;
       pre_pix <= pre_pix;
       proc_in <= proc_in;
       st_ready <= st_ready;
       stencil_0 <= stencil_0;
       stencil_1 <= stencil_1;
       stencil_2 <= stencil_2;
       stencil_3 <= stencil_3;
       stencil_4 <= stencil_4;
       stencil_5 <= stencil_5;
       stencil_6 <= stencil_6;
       stencil_7 <= stencil_7;
       stencil_8 <= stencil_8;
   end
   else if(step) begin
       RAM_w <= n34;
       RAM_x <= n41;
       RAM_y <= n50;
       arg_0_TDATA <= n228;
       arg_0_TVALID <= n239;
       arg_1_TREADY <= n252;
       cur_pix <= n257;
       gbit <= n261;
       pre_pix <= n264;
       proc_in <= n267;
       st_ready <= n270;
       stencil_0 <= n276;
       stencil_1 <= n282;
       stencil_2 <= n288;
       stencil_3 <= n294;
       stencil_4 <= n300;
       stencil_5 <= n306;
       stencil_6 <= n312;
       stencil_7 <= n318;
       stencil_8 <= n404;
       RAM_0 [ RAM_0_addr0 ] <= RAM_0_data0;
       RAM_1 [ RAM_1_addr0 ] <= RAM_1_data0;
       RAM_2 [ RAM_2_addr0 ] <= RAM_2_data0;
       RAM_3 [ RAM_3_addr0 ] <= RAM_3_data0;
       RAM_4 [ RAM_4_addr0 ] <= RAM_4_data0;
       RAM_5 [ RAM_5_addr0 ] <= RAM_5_data0;
       RAM_6 [ RAM_6_addr0 ] <= RAM_6_data0;
       RAM_7 [ RAM_7_addr0 ] <= RAM_7_data0;
   end
end
endmodule
