module riscv(
pc,
x0,
x1,
x10,
x11,
x12,
x13,
x14,
x15,
x16,
x17,
x18,
x19,
x2,
x20,
x21,
x22,
x23,
x24,
x25,
x26,
x27,
x28,
x29,
x3,
x30,
x31,
x4,
x5,
x6,
x7,
x8,
x9,
clk,rst,
step,

// outside memory
mem_raddr0,
mem_rdata0,
mem_raddr1,
mem_rdata1,
mem_raddr2,
mem_rdata2,

mem_wen0,
mem_waddr0,
mem_wdata0
);

output [31:0] mem_raddr0;
output [31:0] mem_raddr1;
output [31:0] mem_raddr2;

input  [31:0] mem_rdata0;
input  [31:0] mem_rdata1;
input  [31:0] mem_rdata2;

output        mem_wen0;
output [31:0] mem_waddr0;
output [31:0] mem_wdata0;


input clk;
input rst;
input step;
output     [31:0] pc;
output     [31:0] x0;
output     [31:0] x1;
output     [31:0] x10;
output     [31:0] x11;
output     [31:0] x12;
output     [31:0] x13;
output     [31:0] x14;
output     [31:0] x15;
output     [31:0] x16;
output     [31:0] x17;
output     [31:0] x18;
output     [31:0] x19;
output     [31:0] x2;
output     [31:0] x20;
output     [31:0] x21;
output     [31:0] x22;
output     [31:0] x23;
output     [31:0] x24;
output     [31:0] x25;
output     [31:0] x26;
output     [31:0] x27;
output     [31:0] x28;
output     [31:0] x29;
output     [31:0] x3;
output     [31:0] x30;
output     [31:0] x31;
output     [31:0] x4;
output     [31:0] x5;
output     [31:0] x6;
output     [31:0] x7;
output     [31:0] x8;
output     [31:0] x9;
reg     [31:0] pc;
reg     [31:0] x0;
reg     [31:0] x1;
reg     [31:0] x10;
reg     [31:0] x11;
reg     [31:0] x12;
reg     [31:0] x13;
reg     [31:0] x14;
reg     [31:0] x15;
reg     [31:0] x16;
reg     [31:0] x17;
reg     [31:0] x18;
reg     [31:0] x19;
reg     [31:0] x2;
reg     [31:0] x20;
reg     [31:0] x21;
reg     [31:0] x22;
reg     [31:0] x23;
reg     [31:0] x24;
reg     [31:0] x25;
reg     [31:0] x26;
reg     [31:0] x27;
reg     [31:0] x28;
reg     [31:0] x29;
reg     [31:0] x3;
reg     [31:0] x30;
reg     [31:0] x31;
reg     [31:0] x4;
reg     [31:0] x5;
reg     [31:0] x6;
reg     [31:0] x7;
reg     [31:0] x8;
reg     [31:0] x9;
wire     [29:0] n0;
wire     [31:0] n1;
wire     [31:0] n2;
wire      [6:0] n3;
wire            n4;
wire      [2:0] n5;
wire            n6;
wire            n7;
wire      [4:0] n8;
wire            n9;
wire            n10;
wire            n11;
wire            n12;
wire            n13;
wire            n14;
wire            n15;
wire            n16;
wire            n17;
wire            n18;
wire            n19;
wire            n20;
wire            n21;
wire            n22;
wire            n23;
wire            n24;
wire            n25;
wire            n26;
wire            n27;
wire            n28;
wire            n29;
wire            n30;
wire            n31;
wire            n32;
wire            n33;
wire            n34;
wire            n35;
wire            n36;
wire            n37;
wire            n38;
wire            n39;
wire     [31:0] n40;
wire     [31:0] n41;
wire     [31:0] n42;
wire     [31:0] n43;
wire     [31:0] n44;
wire     [31:0] n45;
wire     [31:0] n46;
wire     [31:0] n47;
wire     [31:0] n48;
wire     [31:0] n49;
wire     [31:0] n50;
wire     [31:0] n51;
wire     [31:0] n52;
wire     [31:0] n53;
wire     [31:0] n54;
wire     [31:0] n55;
wire     [31:0] n56;
wire     [31:0] n57;
wire     [31:0] n58;
wire     [31:0] n59;
wire     [31:0] n60;
wire     [31:0] n61;
wire     [31:0] n62;
wire     [31:0] n63;
wire     [31:0] n64;
wire     [31:0] n65;
wire     [31:0] n66;
wire     [31:0] n67;
wire     [31:0] n68;
wire     [31:0] n69;
wire     [31:0] n70;
wire     [11:0] n71;
wire     [31:0] n72;
wire     [31:0] n73;
wire     [31:0] n74;
wire            n75;
wire            n76;
wire      [7:0] n77;
wire            n78;
wire      [9:0] n79;
wire     [10:0] n80;
wire     [11:0] n81;
wire     [19:0] n82;
wire     [20:0] n83;
wire     [31:0] n84;
wire     [31:0] n85;
wire            n86;
wire            n87;
wire            n88;
wire      [4:0] n89;
wire            n90;
wire            n91;
wire            n92;
wire            n93;
wire            n94;
wire            n95;
wire            n96;
wire            n97;
wire            n98;
wire            n99;
wire            n100;
wire            n101;
wire            n102;
wire            n103;
wire            n104;
wire            n105;
wire            n106;
wire            n107;
wire            n108;
wire            n109;
wire            n110;
wire            n111;
wire            n112;
wire            n113;
wire            n114;
wire            n115;
wire            n116;
wire            n117;
wire            n118;
wire            n119;
wire            n120;
wire     [31:0] n121;
wire     [31:0] n122;
wire     [31:0] n123;
wire     [31:0] n124;
wire     [31:0] n125;
wire     [31:0] n126;
wire     [31:0] n127;
wire     [31:0] n128;
wire     [31:0] n129;
wire     [31:0] n130;
wire     [31:0] n131;
wire     [31:0] n132;
wire     [31:0] n133;
wire     [31:0] n134;
wire     [31:0] n135;
wire     [31:0] n136;
wire     [31:0] n137;
wire     [31:0] n138;
wire     [31:0] n139;
wire     [31:0] n140;
wire     [31:0] n141;
wire     [31:0] n142;
wire     [31:0] n143;
wire     [31:0] n144;
wire     [31:0] n145;
wire     [31:0] n146;
wire     [31:0] n147;
wire     [31:0] n148;
wire     [31:0] n149;
wire     [31:0] n150;
wire     [31:0] n151;
wire            n152;
wire            n153;
wire      [5:0] n154;
wire      [3:0] n155;
wire      [4:0] n156;
wire     [10:0] n157;
wire     [11:0] n158;
wire     [12:0] n159;
wire     [31:0] n160;
wire     [31:0] n161;
wire     [31:0] n162;
wire     [31:0] n163;
wire            n164;
wire            n165;
wire            n166;
wire     [31:0] n167;
wire            n168;
wire            n169;
wire            n170;
wire     [31:0] n171;
wire            n172;
wire            n173;
wire            n174;
wire     [31:0] n175;
wire            n176;
wire            n177;
wire            n178;
wire     [31:0] n179;
wire            n180;
wire            n181;
wire     [31:0] n182;
wire            n183;
wire            n184;
wire      [6:0] n185;
wire            n186;
wire            n187;
wire            n188;
wire            n189;
wire            n190;
wire            n191;
wire            n192;
wire            n193;
wire            n194;
wire            n195;
wire            n196;
wire            n197;
wire            n198;
wire            n199;
wire            n200;
wire            n201;
wire            n202;
wire            n203;
wire            n204;
wire            n205;
wire            n206;
wire            n207;
wire            n208;
wire            n209;
wire            n210;
wire            n211;
wire            n212;
wire            n213;
wire            n214;
wire            n215;
wire            n216;
wire            n217;
wire            n218;
wire            n219;
wire            n220;
wire            n221;
wire            n222;
wire            n223;
wire            n224;
wire            n225;
wire            n226;
wire            n227;
wire            n228;
wire            n229;
wire            n230;
wire            n231;
wire            n232;
wire            n233;
wire            n234;
wire            n235;
wire            n236;
wire            n237;
wire            n238;
wire            n239;
wire            n240;
wire            n241;
wire            n242;
wire            n243;
wire            n244;
wire            n245;
wire            n246;
wire            n247;
wire            n248;
wire            n249;
wire            n250;
wire            n251;
wire            n252;
wire            n253;
wire            n254;
wire            n255;
wire            n256;
wire            n257;
wire            n258;
wire     [31:0] n259;
wire     [31:0] n260;
wire     [31:0] n261;
wire     [31:0] n262;
wire     [31:0] n263;
wire     [31:0] n264;
wire     [31:0] n265;
wire     [31:0] n266;
wire     [31:0] n267;
wire            n268;
wire            n269;
wire            n270;
wire            n271;
wire            n272;
wire            n273;
wire            n274;
wire            n275;
wire            n276;
wire            n277;
wire            n278;
wire            n279;
wire            n280;
wire            n281;
wire            n282;
wire            n283;
wire            n284;
wire            n285;
wire            n286;
wire            n287;
wire            n288;
wire            n289;
wire            n290;
wire            n291;
wire            n292;
wire            n293;
wire            n294;
wire     [31:0] n295;
wire      [4:0] n296;
wire            n297;
wire      [4:0] n298;
wire     [31:0] n299;
wire     [31:0] n300;
wire     [31:0] n301;
wire     [31:0] n302;
wire     [31:0] n303;
wire     [31:0] n304;
wire     [31:0] n305;
wire     [31:0] n306;
wire     [31:0] n307;
wire     [31:0] n308;
wire     [31:0] n309;
wire     [31:0] n310;
wire     [31:0] n311;
wire     [31:0] n312;
wire     [31:0] n313;
wire     [31:0] n314;
wire     [31:0] n315;
wire     [31:0] n316;
wire     [31:0] n317;
wire     [31:0] n318;
wire     [31:0] n319;
wire     [31:0] n320;
wire     [31:0] n321;
wire     [31:0] n322;
wire     [31:0] n323;
wire     [31:0] n324;
wire     [31:0] n325;
wire     [31:0] n326;
wire     [31:0] n327;
wire     [31:0] n328;
wire     [31:0] n329;
wire     [31:0] n330;
wire     [31:0] n331;
wire     [31:0] n332;
wire     [31:0] n333;
wire     [31:0] n334;
wire            n335;
wire     [31:0] n336;
wire     [31:0] n337;
wire            n338;
wire     [31:0] n339;
wire     [31:0] n340;
wire     [31:0] n341;
wire     [31:0] n342;
wire            n343;
wire     [31:0] n344;
wire     [19:0] n345;
wire     [31:0] n346;
wire     [31:0] n347;
wire     [31:0] n348;
wire     [31:0] n349;
wire      [1:0] n350;
wire            n351;
wire     [29:0] n352;
wire     [31:0] n353;
wire     [31:0] n354;
wire     [15:0] n355;
wire     [31:0] n356;
wire            n357;
wire      [7:0] n358;
wire     [31:0] n359;
wire            n360;
wire     [15:0] n361;
wire     [31:0] n362;
wire            n363;
wire      [7:0] n364;
wire     [31:0] n365;
wire     [31:0] n366;
wire     [31:0] n367;
wire     [31:0] n368;
wire     [31:0] n369;
wire     [31:0] n370;
wire     [31:0] n371;
wire      [7:0] n372;
wire     [31:0] n373;
wire      [7:0] n374;
wire     [31:0] n375;
wire     [31:0] n376;
wire     [31:0] n377;
wire     [31:0] n378;
wire     [31:0] n379;
wire     [31:0] n380;
wire     [31:0] n381;
wire     [31:0] n382;
wire     [31:0] n383;
wire     [31:0] n384;
wire     [31:0] n385;
wire     [31:0] n386;
wire     [31:0] n387;
wire     [31:0] n388;
wire     [31:0] n389;
wire     [31:0] n390;
wire     [31:0] n391;
wire     [31:0] n392;
wire     [31:0] n393;
wire     [31:0] n394;
wire     [31:0] n395;
wire     [31:0] n396;
wire     [31:0] n397;
wire     [31:0] n398;
wire     [31:0] n399;
wire     [31:0] n400;
wire     [31:0] n401;
wire     [31:0] n402;
wire     [31:0] n403;
wire     [31:0] n404;
wire     [31:0] n405;
wire     [31:0] n406;
wire     [31:0] n407;
wire     [31:0] n408;
wire     [31:0] n409;
wire     [31:0] n410;
wire     [31:0] n411;
wire     [31:0] n412;
wire     [31:0] n413;
wire     [31:0] n414;
wire     [31:0] n415;
wire     [31:0] n416;
wire     [31:0] n417;
wire     [31:0] n418;
wire     [31:0] n419;
wire     [31:0] n420;
wire     [31:0] n421;
wire     [31:0] n422;
wire     [31:0] n423;
wire            n424;
wire     [31:0] n425;
wire     [31:0] n426;
wire     [31:0] n427;
wire     [31:0] n428;
wire     [31:0] n429;
wire     [31:0] n430;
wire     [31:0] n431;
wire     [31:0] n432;
wire     [31:0] n433;
wire     [31:0] n434;
wire     [31:0] n435;
wire     [31:0] n436;
wire     [31:0] n437;
wire     [31:0] n438;
wire     [31:0] n439;
wire     [31:0] n440;
wire     [31:0] n441;
wire     [31:0] n442;
wire     [31:0] n443;
wire     [31:0] n444;
wire     [31:0] n445;
wire     [31:0] n446;
wire     [31:0] n447;
wire     [31:0] n448;
wire     [31:0] n449;
wire     [31:0] n450;
wire     [31:0] n451;
wire     [31:0] n452;
wire     [31:0] n453;
wire     [31:0] n454;
wire     [31:0] n455;
wire     [31:0] n456;
wire     [31:0] n457;
wire     [31:0] n458;
wire     [31:0] n459;
wire     [31:0] n460;
wire     [31:0] n461;
wire     [31:0] n462;
wire     [31:0] n463;
wire     [31:0] n464;
wire     [31:0] n465;
wire     [31:0] n466;
wire     [31:0] n467;
wire     [31:0] n468;
wire     [31:0] n469;
wire     [31:0] n470;
wire     [31:0] n471;
wire     [31:0] n472;
wire     [31:0] n473;
wire     [31:0] n474;
wire     [31:0] n475;
wire     [31:0] n476;
wire     [31:0] n477;
wire     [31:0] n478;
wire     [31:0] n479;
wire            n480;
wire     [31:0] n481;
wire     [31:0] n482;
wire     [31:0] n483;
wire     [31:0] n484;
wire     [31:0] n485;
wire     [31:0] n486;
wire     [31:0] n487;
wire     [31:0] n488;
wire     [31:0] n489;
wire     [31:0] n490;
wire     [31:0] n491;
wire     [31:0] n492;
wire     [31:0] n493;
wire     [31:0] n494;
wire     [31:0] n495;
wire     [31:0] n496;
wire     [31:0] n497;
wire     [31:0] n498;
wire     [31:0] n499;
wire     [31:0] n500;
wire     [31:0] n501;
wire     [31:0] n502;
wire     [31:0] n503;
wire     [31:0] n504;
wire     [31:0] n505;
wire     [31:0] n506;
wire     [31:0] n507;
wire     [31:0] n508;
wire     [31:0] n509;
wire     [31:0] n510;
wire     [31:0] n511;
wire     [31:0] n512;
wire     [31:0] n513;
wire     [31:0] n514;
wire     [31:0] n515;
wire     [31:0] n516;
wire     [31:0] n517;
wire     [31:0] n518;
wire     [31:0] n519;
wire     [31:0] n520;
wire     [31:0] n521;
wire     [31:0] n522;
wire     [31:0] n523;
wire     [31:0] n524;
wire     [31:0] n525;
wire     [31:0] n526;
wire     [31:0] n527;
wire     [31:0] n528;
wire     [31:0] n529;
wire     [31:0] n530;
wire     [31:0] n531;
wire     [31:0] n532;
wire     [31:0] n533;
wire     [31:0] n534;
wire            n535;
wire     [31:0] n536;
wire     [31:0] n537;
wire     [31:0] n538;
wire     [31:0] n539;
wire     [31:0] n540;
wire     [31:0] n541;
wire     [31:0] n542;
wire     [31:0] n543;
wire     [31:0] n544;
wire     [31:0] n545;
wire     [31:0] n546;
wire     [31:0] n547;
wire     [31:0] n548;
wire     [31:0] n549;
wire     [31:0] n550;
wire     [31:0] n551;
wire            n552;
wire     [31:0] n553;
wire     [31:0] n554;
wire     [31:0] n555;
wire     [31:0] n556;
wire     [31:0] n557;
wire     [31:0] n558;
wire     [31:0] n559;
wire     [31:0] n560;
wire     [31:0] n561;
wire     [31:0] n562;
wire     [31:0] n563;
wire     [31:0] n564;
wire     [31:0] n565;
wire     [31:0] n566;
wire     [31:0] n567;
wire     [31:0] n568;
wire     [31:0] n569;
wire     [31:0] n570;
wire     [31:0] n571;
wire     [31:0] n572;
wire     [31:0] n573;
wire     [31:0] n574;
wire     [31:0] n575;
wire     [31:0] n576;
wire     [31:0] n577;
wire     [31:0] n578;
wire     [31:0] n579;
wire     [31:0] n580;
wire     [31:0] n581;
wire     [31:0] n582;
wire     [31:0] n583;
wire     [31:0] n584;
wire     [31:0] n585;
wire     [31:0] n586;
wire     [31:0] n587;
wire     [31:0] n588;
wire     [31:0] n589;
wire     [31:0] n590;
wire     [31:0] n591;
wire            n592;
wire     [31:0] n593;
wire     [31:0] n594;
wire     [31:0] n595;
wire     [31:0] n596;
wire     [31:0] n597;
wire     [31:0] n598;
wire     [31:0] n599;
wire     [31:0] n600;
wire     [31:0] n601;
wire     [31:0] n602;
wire     [31:0] n603;
wire     [31:0] n604;
wire     [31:0] n605;
wire     [31:0] n606;
wire     [31:0] n607;
wire     [31:0] n608;
wire     [31:0] n609;
wire     [31:0] n610;
wire            n611;
wire     [31:0] n612;
wire     [31:0] n613;
wire     [31:0] n614;
wire     [31:0] n615;
wire     [31:0] n616;
wire     [31:0] n617;
wire     [31:0] n618;
wire     [31:0] n619;
wire     [31:0] n620;
wire     [31:0] n621;
wire     [31:0] n622;
wire     [31:0] n623;
wire     [31:0] n624;
wire     [31:0] n625;
wire     [31:0] n626;
wire     [31:0] n627;
wire     [31:0] n628;
wire     [31:0] n629;
wire     [31:0] n630;
wire     [31:0] n631;
wire     [31:0] n632;
wire     [31:0] n633;
wire     [31:0] n634;
wire     [31:0] n635;
wire     [31:0] n636;
wire     [31:0] n637;
wire     [31:0] n638;
wire     [31:0] n639;
wire     [31:0] n640;
wire     [31:0] n641;
wire     [31:0] n642;
wire     [31:0] n643;
wire     [31:0] n644;
wire     [31:0] n645;
wire     [31:0] n646;
wire     [31:0] n647;
wire     [31:0] n648;
wire     [31:0] n649;
wire            n650;
wire     [31:0] n651;
wire     [31:0] n652;
wire     [31:0] n653;
wire     [31:0] n654;
wire     [31:0] n655;
wire     [31:0] n656;
wire     [31:0] n657;
wire     [31:0] n658;
wire     [31:0] n659;
wire     [31:0] n660;
wire     [31:0] n661;
wire     [31:0] n662;
wire     [31:0] n663;
wire     [31:0] n664;
wire     [31:0] n665;
wire     [31:0] n666;
wire     [31:0] n667;
wire     [31:0] n668;
wire     [31:0] n669;
wire     [31:0] n670;
wire     [31:0] n671;
wire     [31:0] n672;
wire     [31:0] n673;
wire     [31:0] n674;
wire     [31:0] n675;
wire     [31:0] n676;
wire     [31:0] n677;
wire     [31:0] n678;
wire     [31:0] n679;
wire     [31:0] n680;
wire     [31:0] n681;
wire     [31:0] n682;
wire     [31:0] n683;
wire     [31:0] n684;
wire     [31:0] n685;
wire     [31:0] n686;
wire     [31:0] n687;
wire     [31:0] n688;
wire     [31:0] n689;
wire     [31:0] n690;
wire     [31:0] n691;
wire     [31:0] n692;
wire     [31:0] n693;
wire     [31:0] n694;
wire     [31:0] n695;
wire     [31:0] n696;
wire     [31:0] n697;
wire     [31:0] n698;
wire     [31:0] n699;
wire     [31:0] n700;
wire     [31:0] n701;
wire     [31:0] n702;
wire     [31:0] n703;
wire     [31:0] n704;
wire            n705;
wire     [31:0] n706;
wire     [31:0] n707;
wire     [31:0] n708;
wire     [31:0] n709;
wire     [31:0] n710;
wire     [31:0] n711;
wire     [31:0] n712;
wire     [31:0] n713;
wire     [31:0] n714;
wire     [31:0] n715;
wire     [31:0] n716;
wire     [31:0] n717;
wire     [31:0] n718;
wire     [31:0] n719;
wire     [31:0] n720;
wire     [31:0] n721;
wire     [31:0] n722;
wire     [31:0] n723;
wire     [31:0] n724;
wire     [31:0] n725;
wire     [31:0] n726;
wire     [31:0] n727;
wire     [31:0] n728;
wire     [31:0] n729;
wire     [31:0] n730;
wire     [31:0] n731;
wire     [31:0] n732;
wire     [31:0] n733;
wire     [31:0] n734;
wire     [31:0] n735;
wire     [31:0] n736;
wire     [31:0] n737;
wire     [31:0] n738;
wire     [31:0] n739;
wire     [31:0] n740;
wire     [31:0] n741;
wire     [31:0] n742;
wire     [31:0] n743;
wire     [31:0] n744;
wire     [31:0] n745;
wire     [31:0] n746;
wire     [31:0] n747;
wire     [31:0] n748;
wire     [31:0] n749;
wire     [31:0] n750;
wire     [31:0] n751;
wire     [31:0] n752;
wire     [31:0] n753;
wire     [31:0] n754;
wire     [31:0] n755;
wire     [31:0] n756;
wire     [31:0] n757;
wire     [31:0] n758;
wire     [31:0] n759;
wire     [31:0] n760;
wire            n761;
wire     [31:0] n762;
wire     [31:0] n763;
wire     [31:0] n764;
wire     [31:0] n765;
wire     [31:0] n766;
wire     [31:0] n767;
wire     [31:0] n768;
wire     [31:0] n769;
wire     [31:0] n770;
wire     [31:0] n771;
wire     [31:0] n772;
wire     [31:0] n773;
wire     [31:0] n774;
wire     [31:0] n775;
wire     [31:0] n776;
wire     [31:0] n777;
wire     [31:0] n778;
wire     [31:0] n779;
wire     [31:0] n780;
wire     [31:0] n781;
wire     [31:0] n782;
wire     [31:0] n783;
wire     [31:0] n784;
wire     [31:0] n785;
wire     [31:0] n786;
wire     [31:0] n787;
wire     [31:0] n788;
wire     [31:0] n789;
wire     [31:0] n790;
wire     [31:0] n791;
wire     [31:0] n792;
wire     [31:0] n793;
wire     [31:0] n794;
wire     [31:0] n795;
wire     [31:0] n796;
wire     [31:0] n797;
wire     [31:0] n798;
wire     [31:0] n799;
wire     [31:0] n800;
wire     [31:0] n801;
wire     [31:0] n802;
wire     [31:0] n803;
wire     [31:0] n804;
wire     [31:0] n805;
wire     [31:0] n806;
wire     [31:0] n807;
wire     [31:0] n808;
wire     [31:0] n809;
wire     [31:0] n810;
wire     [31:0] n811;
wire     [31:0] n812;
wire     [31:0] n813;
wire     [31:0] n814;
wire     [31:0] n815;
wire            n816;
wire     [31:0] n817;
wire     [31:0] n818;
wire     [31:0] n819;
wire     [31:0] n820;
wire     [31:0] n821;
wire     [31:0] n822;
wire     [31:0] n823;
wire     [31:0] n824;
wire     [31:0] n825;
wire     [31:0] n826;
wire     [31:0] n827;
wire     [31:0] n828;
wire     [31:0] n829;
wire     [31:0] n830;
wire     [31:0] n831;
wire     [31:0] n832;
wire     [31:0] n833;
wire     [31:0] n834;
wire     [31:0] n835;
wire     [31:0] n836;
wire     [31:0] n837;
wire     [31:0] n838;
wire     [31:0] n839;
wire     [31:0] n840;
wire     [31:0] n841;
wire     [31:0] n842;
wire     [31:0] n843;
wire     [31:0] n844;
wire     [31:0] n845;
wire     [31:0] n846;
wire     [31:0] n847;
wire     [31:0] n848;
wire     [31:0] n849;
wire     [31:0] n850;
wire     [31:0] n851;
wire     [31:0] n852;
wire     [31:0] n853;
wire     [31:0] n854;
wire     [31:0] n855;
wire     [31:0] n856;
wire     [31:0] n857;
wire     [31:0] n858;
wire     [31:0] n859;
wire     [31:0] n860;
wire     [31:0] n861;
wire     [31:0] n862;
wire     [31:0] n863;
wire     [31:0] n864;
wire     [31:0] n865;
wire     [31:0] n866;
wire     [31:0] n867;
wire     [31:0] n868;
wire     [31:0] n869;
wire     [31:0] n870;
wire            n871;
wire     [31:0] n872;
wire     [31:0] n873;
wire     [31:0] n874;
wire     [31:0] n875;
wire     [31:0] n876;
wire     [31:0] n877;
wire     [31:0] n878;
wire     [31:0] n879;
wire     [31:0] n880;
wire     [31:0] n881;
wire     [31:0] n882;
wire     [31:0] n883;
wire     [31:0] n884;
wire     [31:0] n885;
wire     [31:0] n886;
wire     [31:0] n887;
wire     [31:0] n888;
wire     [31:0] n889;
wire     [31:0] n890;
wire     [31:0] n891;
wire     [31:0] n892;
wire     [31:0] n893;
wire     [31:0] n894;
wire     [31:0] n895;
wire     [31:0] n896;
wire     [31:0] n897;
wire     [31:0] n898;
wire     [31:0] n899;
wire     [31:0] n900;
wire     [31:0] n901;
wire     [31:0] n902;
wire     [31:0] n903;
wire     [31:0] n904;
wire     [31:0] n905;
wire     [31:0] n906;
wire     [31:0] n907;
wire     [31:0] n908;
wire     [31:0] n909;
wire     [31:0] n910;
wire     [31:0] n911;
wire     [31:0] n912;
wire     [31:0] n913;
wire     [31:0] n914;
wire     [31:0] n915;
wire     [31:0] n916;
wire     [31:0] n917;
wire     [31:0] n918;
wire     [31:0] n919;
wire     [31:0] n920;
wire     [31:0] n921;
wire     [31:0] n922;
wire     [31:0] n923;
wire     [31:0] n924;
wire     [31:0] n925;
wire            n926;
wire     [31:0] n927;
wire     [31:0] n928;
wire     [31:0] n929;
wire     [31:0] n930;
wire     [31:0] n931;
wire     [31:0] n932;
wire     [31:0] n933;
wire     [31:0] n934;
wire     [31:0] n935;
wire     [31:0] n936;
wire     [31:0] n937;
wire     [31:0] n938;
wire     [31:0] n939;
wire     [31:0] n940;
wire     [31:0] n941;
wire     [31:0] n942;
wire     [31:0] n943;
wire     [31:0] n944;
wire     [31:0] n945;
wire     [31:0] n946;
wire     [31:0] n947;
wire     [31:0] n948;
wire     [31:0] n949;
wire     [31:0] n950;
wire     [31:0] n951;
wire     [31:0] n952;
wire     [31:0] n953;
wire     [31:0] n954;
wire     [31:0] n955;
wire     [31:0] n956;
wire     [31:0] n957;
wire     [31:0] n958;
wire     [31:0] n959;
wire     [31:0] n960;
wire     [31:0] n961;
wire     [31:0] n962;
wire     [31:0] n963;
wire     [31:0] n964;
wire     [31:0] n965;
wire     [31:0] n966;
wire     [31:0] n967;
wire     [31:0] n968;
wire     [31:0] n969;
wire     [31:0] n970;
wire     [31:0] n971;
wire     [31:0] n972;
wire     [31:0] n973;
wire     [31:0] n974;
wire     [31:0] n975;
wire     [31:0] n976;
wire     [31:0] n977;
wire     [31:0] n978;
wire     [31:0] n979;
wire     [31:0] n980;
wire            n981;
wire     [31:0] n982;
wire     [31:0] n983;
wire     [31:0] n984;
wire     [31:0] n985;
wire     [31:0] n986;
wire     [31:0] n987;
wire     [31:0] n988;
wire     [31:0] n989;
wire     [31:0] n990;
wire     [31:0] n991;
wire     [31:0] n992;
wire     [31:0] n993;
wire     [31:0] n994;
wire     [31:0] n995;
wire     [31:0] n996;
wire     [31:0] n997;
wire     [31:0] n998;
wire     [31:0] n999;
wire     [31:0] n1000;
wire     [31:0] n1001;
wire     [31:0] n1002;
wire     [31:0] n1003;
wire     [31:0] n1004;
wire     [31:0] n1005;
wire     [31:0] n1006;
wire     [31:0] n1007;
wire     [31:0] n1008;
wire     [31:0] n1009;
wire     [31:0] n1010;
wire     [31:0] n1011;
wire     [31:0] n1012;
wire     [31:0] n1013;
wire     [31:0] n1014;
wire     [31:0] n1015;
wire     [31:0] n1016;
wire     [31:0] n1017;
wire     [31:0] n1018;
wire     [31:0] n1019;
wire     [31:0] n1020;
wire     [31:0] n1021;
wire     [31:0] n1022;
wire     [31:0] n1023;
wire     [31:0] n1024;
wire     [31:0] n1025;
wire     [31:0] n1026;
wire     [31:0] n1027;
wire     [31:0] n1028;
wire     [31:0] n1029;
wire     [31:0] n1030;
wire     [31:0] n1031;
wire     [31:0] n1032;
wire     [31:0] n1033;
wire     [31:0] n1034;
wire     [31:0] n1035;
wire            n1036;
wire     [31:0] n1037;
wire     [31:0] n1038;
wire     [31:0] n1039;
wire     [31:0] n1040;
wire     [31:0] n1041;
wire     [31:0] n1042;
wire     [31:0] n1043;
wire     [31:0] n1044;
wire     [31:0] n1045;
wire     [31:0] n1046;
wire     [31:0] n1047;
wire     [31:0] n1048;
wire     [31:0] n1049;
wire     [31:0] n1050;
wire     [31:0] n1051;
wire     [31:0] n1052;
wire     [31:0] n1053;
wire     [31:0] n1054;
wire     [31:0] n1055;
wire     [31:0] n1056;
wire     [31:0] n1057;
wire     [31:0] n1058;
wire     [31:0] n1059;
wire     [31:0] n1060;
wire     [31:0] n1061;
wire     [31:0] n1062;
wire     [31:0] n1063;
wire     [31:0] n1064;
wire     [31:0] n1065;
wire     [31:0] n1066;
wire     [31:0] n1067;
wire     [31:0] n1068;
wire     [31:0] n1069;
wire     [31:0] n1070;
wire     [31:0] n1071;
wire     [31:0] n1072;
wire     [31:0] n1073;
wire     [31:0] n1074;
wire     [31:0] n1075;
wire     [31:0] n1076;
wire     [31:0] n1077;
wire     [31:0] n1078;
wire     [31:0] n1079;
wire     [31:0] n1080;
wire     [31:0] n1081;
wire     [31:0] n1082;
wire     [31:0] n1083;
wire     [31:0] n1084;
wire     [31:0] n1085;
wire     [31:0] n1086;
wire     [31:0] n1087;
wire     [31:0] n1088;
wire     [31:0] n1089;
wire     [31:0] n1090;
wire            n1091;
wire     [31:0] n1092;
wire     [31:0] n1093;
wire     [31:0] n1094;
wire     [31:0] n1095;
wire     [31:0] n1096;
wire     [31:0] n1097;
wire     [31:0] n1098;
wire     [31:0] n1099;
wire     [31:0] n1100;
wire     [31:0] n1101;
wire     [31:0] n1102;
wire     [31:0] n1103;
wire     [31:0] n1104;
wire     [31:0] n1105;
wire     [31:0] n1106;
wire     [31:0] n1107;
wire     [31:0] n1108;
wire     [31:0] n1109;
wire     [31:0] n1110;
wire     [31:0] n1111;
wire     [31:0] n1112;
wire     [31:0] n1113;
wire     [31:0] n1114;
wire     [31:0] n1115;
wire     [31:0] n1116;
wire     [31:0] n1117;
wire     [31:0] n1118;
wire     [31:0] n1119;
wire     [31:0] n1120;
wire     [31:0] n1121;
wire     [31:0] n1122;
wire     [31:0] n1123;
wire     [31:0] n1124;
wire     [31:0] n1125;
wire     [31:0] n1126;
wire     [31:0] n1127;
wire     [31:0] n1128;
wire     [31:0] n1129;
wire     [31:0] n1130;
wire     [31:0] n1131;
wire     [31:0] n1132;
wire     [31:0] n1133;
wire     [31:0] n1134;
wire     [31:0] n1135;
wire     [31:0] n1136;
wire     [31:0] n1137;
wire     [31:0] n1138;
wire     [31:0] n1139;
wire     [31:0] n1140;
wire     [31:0] n1141;
wire     [31:0] n1142;
wire     [31:0] n1143;
wire     [31:0] n1144;
wire     [31:0] n1145;
wire            n1146;
wire     [31:0] n1147;
wire     [31:0] n1148;
wire     [31:0] n1149;
wire     [31:0] n1150;
wire     [31:0] n1151;
wire     [31:0] n1152;
wire     [31:0] n1153;
wire     [31:0] n1154;
wire     [31:0] n1155;
wire     [31:0] n1156;
wire     [31:0] n1157;
wire     [31:0] n1158;
wire     [31:0] n1159;
wire     [31:0] n1160;
wire     [31:0] n1161;
wire     [31:0] n1162;
wire     [31:0] n1163;
wire     [31:0] n1164;
wire     [31:0] n1165;
wire     [31:0] n1166;
wire     [31:0] n1167;
wire     [31:0] n1168;
wire     [31:0] n1169;
wire     [31:0] n1170;
wire     [31:0] n1171;
wire     [31:0] n1172;
wire     [31:0] n1173;
wire     [31:0] n1174;
wire     [31:0] n1175;
wire     [31:0] n1176;
wire     [31:0] n1177;
wire     [31:0] n1178;
wire     [31:0] n1179;
wire     [31:0] n1180;
wire     [31:0] n1181;
wire     [31:0] n1182;
wire     [31:0] n1183;
wire     [31:0] n1184;
wire     [31:0] n1185;
wire     [31:0] n1186;
wire     [31:0] n1187;
wire     [31:0] n1188;
wire     [31:0] n1189;
wire     [31:0] n1190;
wire     [31:0] n1191;
wire     [31:0] n1192;
wire     [31:0] n1193;
wire     [31:0] n1194;
wire     [31:0] n1195;
wire     [31:0] n1196;
wire     [31:0] n1197;
wire     [31:0] n1198;
wire     [31:0] n1199;
wire     [31:0] n1200;
wire            n1201;
wire     [31:0] n1202;
wire     [31:0] n1203;
wire     [31:0] n1204;
wire     [31:0] n1205;
wire     [31:0] n1206;
wire     [31:0] n1207;
wire     [31:0] n1208;
wire     [31:0] n1209;
wire     [31:0] n1210;
wire     [31:0] n1211;
wire     [31:0] n1212;
wire     [31:0] n1213;
wire     [31:0] n1214;
wire     [31:0] n1215;
wire     [31:0] n1216;
wire     [31:0] n1217;
wire     [31:0] n1218;
wire     [31:0] n1219;
wire     [31:0] n1220;
wire     [31:0] n1221;
wire     [31:0] n1222;
wire     [31:0] n1223;
wire     [31:0] n1224;
wire     [31:0] n1225;
wire     [31:0] n1226;
wire     [31:0] n1227;
wire     [31:0] n1228;
wire     [31:0] n1229;
wire     [31:0] n1230;
wire     [31:0] n1231;
wire     [31:0] n1232;
wire     [31:0] n1233;
wire     [31:0] n1234;
wire     [31:0] n1235;
wire     [31:0] n1236;
wire     [31:0] n1237;
wire     [31:0] n1238;
wire     [31:0] n1239;
wire     [31:0] n1240;
wire     [31:0] n1241;
wire     [31:0] n1242;
wire     [31:0] n1243;
wire     [31:0] n1244;
wire     [31:0] n1245;
wire     [31:0] n1246;
wire     [31:0] n1247;
wire     [31:0] n1248;
wire     [31:0] n1249;
wire     [31:0] n1250;
wire     [31:0] n1251;
wire     [31:0] n1252;
wire     [31:0] n1253;
wire     [31:0] n1254;
wire     [31:0] n1255;
wire            n1256;
wire     [31:0] n1257;
wire     [31:0] n1258;
wire     [31:0] n1259;
wire     [31:0] n1260;
wire     [31:0] n1261;
wire     [31:0] n1262;
wire     [31:0] n1263;
wire     [31:0] n1264;
wire     [31:0] n1265;
wire     [31:0] n1266;
wire     [31:0] n1267;
wire     [31:0] n1268;
wire     [31:0] n1269;
wire     [31:0] n1270;
wire     [31:0] n1271;
wire     [31:0] n1272;
wire     [31:0] n1273;
wire     [31:0] n1274;
wire     [31:0] n1275;
wire     [31:0] n1276;
wire     [31:0] n1277;
wire     [31:0] n1278;
wire     [31:0] n1279;
wire     [31:0] n1280;
wire     [31:0] n1281;
wire     [31:0] n1282;
wire     [31:0] n1283;
wire     [31:0] n1284;
wire     [31:0] n1285;
wire     [31:0] n1286;
wire     [31:0] n1287;
wire     [31:0] n1288;
wire     [31:0] n1289;
wire     [31:0] n1290;
wire     [31:0] n1291;
wire     [31:0] n1292;
wire     [31:0] n1293;
wire     [31:0] n1294;
wire     [31:0] n1295;
wire     [31:0] n1296;
wire     [31:0] n1297;
wire     [31:0] n1298;
wire     [31:0] n1299;
wire     [31:0] n1300;
wire     [31:0] n1301;
wire     [31:0] n1302;
wire     [31:0] n1303;
wire     [31:0] n1304;
wire     [31:0] n1305;
wire     [31:0] n1306;
wire     [31:0] n1307;
wire     [31:0] n1308;
wire     [31:0] n1309;
wire     [31:0] n1310;
wire            n1311;
wire     [31:0] n1312;
wire     [31:0] n1313;
wire     [31:0] n1314;
wire     [31:0] n1315;
wire     [31:0] n1316;
wire     [31:0] n1317;
wire     [31:0] n1318;
wire     [31:0] n1319;
wire     [31:0] n1320;
wire     [31:0] n1321;
wire     [31:0] n1322;
wire     [31:0] n1323;
wire     [31:0] n1324;
wire     [31:0] n1325;
wire     [31:0] n1326;
wire     [31:0] n1327;
wire     [31:0] n1328;
wire     [31:0] n1329;
wire     [31:0] n1330;
wire     [31:0] n1331;
wire     [31:0] n1332;
wire     [31:0] n1333;
wire     [31:0] n1334;
wire     [31:0] n1335;
wire     [31:0] n1336;
wire     [31:0] n1337;
wire     [31:0] n1338;
wire     [31:0] n1339;
wire     [31:0] n1340;
wire     [31:0] n1341;
wire     [31:0] n1342;
wire     [31:0] n1343;
wire     [31:0] n1344;
wire     [31:0] n1345;
wire     [31:0] n1346;
wire     [31:0] n1347;
wire     [31:0] n1348;
wire     [31:0] n1349;
wire     [31:0] n1350;
wire     [31:0] n1351;
wire     [31:0] n1352;
wire     [31:0] n1353;
wire     [31:0] n1354;
wire     [31:0] n1355;
wire     [31:0] n1356;
wire     [31:0] n1357;
wire     [31:0] n1358;
wire     [31:0] n1359;
wire     [31:0] n1360;
wire     [31:0] n1361;
wire     [31:0] n1362;
wire     [31:0] n1363;
wire     [31:0] n1364;
wire     [31:0] n1365;
wire            n1366;
wire     [31:0] n1367;
wire     [31:0] n1368;
wire     [31:0] n1369;
wire     [31:0] n1370;
wire     [31:0] n1371;
wire     [31:0] n1372;
wire     [31:0] n1373;
wire     [31:0] n1374;
wire     [31:0] n1375;
wire     [31:0] n1376;
wire     [31:0] n1377;
wire     [31:0] n1378;
wire     [31:0] n1379;
wire     [31:0] n1380;
wire     [31:0] n1381;
wire     [31:0] n1382;
wire     [31:0] n1383;
wire     [31:0] n1384;
wire     [31:0] n1385;
wire     [31:0] n1386;
wire     [31:0] n1387;
wire     [31:0] n1388;
wire     [31:0] n1389;
wire     [31:0] n1390;
wire     [31:0] n1391;
wire     [31:0] n1392;
wire     [31:0] n1393;
wire     [31:0] n1394;
wire     [31:0] n1395;
wire     [31:0] n1396;
wire     [31:0] n1397;
wire     [31:0] n1398;
wire     [31:0] n1399;
wire     [31:0] n1400;
wire     [31:0] n1401;
wire     [31:0] n1402;
wire     [31:0] n1403;
wire     [31:0] n1404;
wire     [31:0] n1405;
wire     [31:0] n1406;
wire     [31:0] n1407;
wire     [31:0] n1408;
wire     [31:0] n1409;
wire     [31:0] n1410;
wire     [31:0] n1411;
wire     [31:0] n1412;
wire     [31:0] n1413;
wire     [31:0] n1414;
wire     [31:0] n1415;
wire     [31:0] n1416;
wire     [31:0] n1417;
wire     [31:0] n1418;
wire     [31:0] n1419;
wire     [31:0] n1420;
wire            n1421;
wire     [31:0] n1422;
wire     [31:0] n1423;
wire     [31:0] n1424;
wire     [31:0] n1425;
wire     [31:0] n1426;
wire     [31:0] n1427;
wire     [31:0] n1428;
wire     [31:0] n1429;
wire     [31:0] n1430;
wire     [31:0] n1431;
wire     [31:0] n1432;
wire     [31:0] n1433;
wire     [31:0] n1434;
wire     [31:0] n1435;
wire     [31:0] n1436;
wire     [31:0] n1437;
wire     [31:0] n1438;
wire     [31:0] n1439;
wire     [31:0] n1440;
wire     [31:0] n1441;
wire     [31:0] n1442;
wire     [31:0] n1443;
wire     [31:0] n1444;
wire     [31:0] n1445;
wire     [31:0] n1446;
wire     [31:0] n1447;
wire     [31:0] n1448;
wire     [31:0] n1449;
wire     [31:0] n1450;
wire     [31:0] n1451;
wire     [31:0] n1452;
wire     [31:0] n1453;
wire     [31:0] n1454;
wire     [31:0] n1455;
wire     [31:0] n1456;
wire     [31:0] n1457;
wire     [31:0] n1458;
wire     [31:0] n1459;
wire     [31:0] n1460;
wire     [31:0] n1461;
wire     [31:0] n1462;
wire     [31:0] n1463;
wire     [31:0] n1464;
wire     [31:0] n1465;
wire     [31:0] n1466;
wire     [31:0] n1467;
wire     [31:0] n1468;
wire     [31:0] n1469;
wire     [31:0] n1470;
wire     [31:0] n1471;
wire     [31:0] n1472;
wire     [31:0] n1473;
wire     [31:0] n1474;
wire     [31:0] n1475;
wire            n1476;
wire     [31:0] n1477;
wire     [31:0] n1478;
wire     [31:0] n1479;
wire     [31:0] n1480;
wire     [31:0] n1481;
wire     [31:0] n1482;
wire     [31:0] n1483;
wire     [31:0] n1484;
wire     [31:0] n1485;
wire     [31:0] n1486;
wire     [31:0] n1487;
wire     [31:0] n1488;
wire     [31:0] n1489;
wire     [31:0] n1490;
wire     [31:0] n1491;
wire     [31:0] n1492;
wire     [31:0] n1493;
wire     [31:0] n1494;
wire     [31:0] n1495;
wire     [31:0] n1496;
wire     [31:0] n1497;
wire     [31:0] n1498;
wire     [31:0] n1499;
wire     [31:0] n1500;
wire     [31:0] n1501;
wire     [31:0] n1502;
wire     [31:0] n1503;
wire     [31:0] n1504;
wire     [31:0] n1505;
wire     [31:0] n1506;
wire     [31:0] n1507;
wire     [31:0] n1508;
wire     [31:0] n1509;
wire     [31:0] n1510;
wire     [31:0] n1511;
wire     [31:0] n1512;
wire     [31:0] n1513;
wire     [31:0] n1514;
wire     [31:0] n1515;
wire     [31:0] n1516;
wire     [31:0] n1517;
wire     [31:0] n1518;
wire     [31:0] n1519;
wire     [31:0] n1520;
wire     [31:0] n1521;
wire     [31:0] n1522;
wire     [31:0] n1523;
wire     [31:0] n1524;
wire     [31:0] n1525;
wire     [31:0] n1526;
wire     [31:0] n1527;
wire     [31:0] n1528;
wire     [31:0] n1529;
wire     [31:0] n1530;
wire            n1531;
wire     [31:0] n1532;
wire     [31:0] n1533;
wire     [31:0] n1534;
wire     [31:0] n1535;
wire     [31:0] n1536;
wire     [31:0] n1537;
wire     [31:0] n1538;
wire     [31:0] n1539;
wire     [31:0] n1540;
wire     [31:0] n1541;
wire     [31:0] n1542;
wire     [31:0] n1543;
wire     [31:0] n1544;
wire     [31:0] n1545;
wire     [31:0] n1546;
wire     [31:0] n1547;
wire     [31:0] n1548;
wire     [31:0] n1549;
wire     [31:0] n1550;
wire     [31:0] n1551;
wire     [31:0] n1552;
wire     [31:0] n1553;
wire     [31:0] n1554;
wire     [31:0] n1555;
wire     [31:0] n1556;
wire     [31:0] n1557;
wire     [31:0] n1558;
wire     [31:0] n1559;
wire     [31:0] n1560;
wire     [31:0] n1561;
wire     [31:0] n1562;
wire     [31:0] n1563;
wire     [31:0] n1564;
wire     [31:0] n1565;
wire     [31:0] n1566;
wire     [31:0] n1567;
wire     [31:0] n1568;
wire     [31:0] n1569;
wire     [31:0] n1570;
wire     [31:0] n1571;
wire     [31:0] n1572;
wire     [31:0] n1573;
wire     [31:0] n1574;
wire     [31:0] n1575;
wire     [31:0] n1576;
wire     [31:0] n1577;
wire     [31:0] n1578;
wire     [31:0] n1579;
wire     [31:0] n1580;
wire     [31:0] n1581;
wire     [31:0] n1582;
wire     [31:0] n1583;
wire     [31:0] n1584;
wire     [31:0] n1585;
wire            n1586;
wire     [31:0] n1587;
wire     [31:0] n1588;
wire     [31:0] n1589;
wire     [31:0] n1590;
wire     [31:0] n1591;
wire     [31:0] n1592;
wire     [31:0] n1593;
wire     [31:0] n1594;
wire     [31:0] n1595;
wire     [31:0] n1596;
wire     [31:0] n1597;
wire     [31:0] n1598;
wire     [31:0] n1599;
wire     [31:0] n1600;
wire     [31:0] n1601;
wire     [31:0] n1602;
wire     [31:0] n1603;
wire     [31:0] n1604;
wire     [31:0] n1605;
wire     [31:0] n1606;
wire     [31:0] n1607;
wire     [31:0] n1608;
wire     [31:0] n1609;
wire     [31:0] n1610;
wire     [31:0] n1611;
wire     [31:0] n1612;
wire     [31:0] n1613;
wire     [31:0] n1614;
wire     [31:0] n1615;
wire     [31:0] n1616;
wire     [31:0] n1617;
wire     [31:0] n1618;
wire     [31:0] n1619;
wire     [31:0] n1620;
wire     [31:0] n1621;
wire     [31:0] n1622;
wire     [31:0] n1623;
wire     [31:0] n1624;
wire     [31:0] n1625;
wire     [31:0] n1626;
wire     [31:0] n1627;
wire     [31:0] n1628;
wire     [31:0] n1629;
wire     [31:0] n1630;
wire     [31:0] n1631;
wire     [31:0] n1632;
wire     [31:0] n1633;
wire     [31:0] n1634;
wire     [31:0] n1635;
wire     [31:0] n1636;
wire     [31:0] n1637;
wire     [31:0] n1638;
wire     [31:0] n1639;
wire     [31:0] n1640;
wire            n1641;
wire     [31:0] n1642;
wire     [31:0] n1643;
wire     [31:0] n1644;
wire     [31:0] n1645;
wire     [31:0] n1646;
wire     [31:0] n1647;
wire     [31:0] n1648;
wire     [31:0] n1649;
wire     [31:0] n1650;
wire     [31:0] n1651;
wire     [31:0] n1652;
wire     [31:0] n1653;
wire     [31:0] n1654;
wire     [31:0] n1655;
wire     [31:0] n1656;
wire     [31:0] n1657;
wire     [31:0] n1658;
wire     [31:0] n1659;
wire     [31:0] n1660;
wire     [31:0] n1661;
wire     [31:0] n1662;
wire     [31:0] n1663;
wire     [31:0] n1664;
wire     [31:0] n1665;
wire     [31:0] n1666;
wire     [31:0] n1667;
wire     [31:0] n1668;
wire     [31:0] n1669;
wire     [31:0] n1670;
wire     [31:0] n1671;
wire     [31:0] n1672;
wire     [31:0] n1673;
wire     [31:0] n1674;
wire     [31:0] n1675;
wire     [31:0] n1676;
wire     [31:0] n1677;
wire     [31:0] n1678;
wire     [31:0] n1679;
wire     [31:0] n1680;
wire     [31:0] n1681;
wire     [31:0] n1682;
wire     [31:0] n1683;
wire     [31:0] n1684;
wire     [31:0] n1685;
wire     [31:0] n1686;
wire     [31:0] n1687;
wire     [31:0] n1688;
wire     [31:0] n1689;
wire     [31:0] n1690;
wire     [31:0] n1691;
wire     [31:0] n1692;
wire     [31:0] n1693;
wire     [31:0] n1694;
wire     [31:0] n1695;
wire            n1696;
wire     [31:0] n1697;
wire     [31:0] n1698;
wire     [31:0] n1699;
wire     [31:0] n1700;
wire     [31:0] n1701;
wire     [31:0] n1702;
wire     [31:0] n1703;
wire     [31:0] n1704;
wire     [31:0] n1705;
wire     [31:0] n1706;
wire     [31:0] n1707;
wire     [31:0] n1708;
wire     [31:0] n1709;
wire     [31:0] n1710;
wire     [31:0] n1711;
wire     [31:0] n1712;
wire     [31:0] n1713;
wire     [31:0] n1714;
wire     [31:0] n1715;
wire     [31:0] n1716;
wire     [31:0] n1717;
wire     [31:0] n1718;
wire     [31:0] n1719;
wire     [31:0] n1720;
wire     [31:0] n1721;
wire     [31:0] n1722;
wire     [31:0] n1723;
wire     [31:0] n1724;
wire     [31:0] n1725;
wire     [31:0] n1726;
wire     [31:0] n1727;
wire     [31:0] n1728;
wire     [31:0] n1729;
wire     [31:0] n1730;
wire     [31:0] n1731;
wire     [31:0] n1732;
wire     [31:0] n1733;
wire     [31:0] n1734;
wire     [31:0] n1735;
wire     [31:0] n1736;
wire     [31:0] n1737;
wire     [31:0] n1738;
wire     [31:0] n1739;
wire     [31:0] n1740;
wire     [31:0] n1741;
wire     [31:0] n1742;
wire     [31:0] n1743;
wire     [31:0] n1744;
wire     [31:0] n1745;
wire     [31:0] n1746;
wire     [31:0] n1747;
wire     [31:0] n1748;
wire     [31:0] n1749;
wire     [31:0] n1750;
wire            n1751;
wire     [31:0] n1752;
wire     [31:0] n1753;
wire     [31:0] n1754;
wire     [31:0] n1755;
wire     [31:0] n1756;
wire     [31:0] n1757;
wire     [31:0] n1758;
wire     [31:0] n1759;
wire     [31:0] n1760;
wire     [31:0] n1761;
wire     [31:0] n1762;
wire     [31:0] n1763;
wire     [31:0] n1764;
wire     [31:0] n1765;
wire     [31:0] n1766;
wire     [31:0] n1767;
wire     [31:0] n1768;
wire     [31:0] n1769;
wire     [31:0] n1770;
wire     [31:0] n1771;
wire     [31:0] n1772;
wire     [31:0] n1773;
wire     [31:0] n1774;
wire     [31:0] n1775;
wire     [31:0] n1776;
wire     [31:0] n1777;
wire     [31:0] n1778;
wire     [31:0] n1779;
wire     [31:0] n1780;
wire     [31:0] n1781;
wire     [31:0] n1782;
wire     [31:0] n1783;
wire     [31:0] n1784;
wire     [31:0] n1785;
wire     [31:0] n1786;
wire     [31:0] n1787;
wire     [31:0] n1788;
wire     [31:0] n1789;
wire     [31:0] n1790;
wire     [31:0] n1791;
wire     [31:0] n1792;
wire     [31:0] n1793;
wire     [31:0] n1794;
wire     [31:0] n1795;
wire     [31:0] n1796;
wire     [31:0] n1797;
wire     [31:0] n1798;
wire     [31:0] n1799;
wire     [31:0] n1800;
wire     [31:0] n1801;
wire     [31:0] n1802;
wire     [31:0] n1803;
wire     [31:0] n1804;
wire     [31:0] n1805;
wire            n1806;
wire     [31:0] n1807;
wire     [31:0] n1808;
wire     [31:0] n1809;
wire     [31:0] n1810;
wire     [31:0] n1811;
wire     [31:0] n1812;
wire     [31:0] n1813;
wire     [31:0] n1814;
wire     [31:0] n1815;
wire     [31:0] n1816;
wire     [31:0] n1817;
wire     [31:0] n1818;
wire     [31:0] n1819;
wire     [31:0] n1820;
wire     [31:0] n1821;
wire     [31:0] n1822;
wire     [31:0] n1823;
wire     [31:0] n1824;
wire     [31:0] n1825;
wire     [31:0] n1826;
wire     [31:0] n1827;
wire     [31:0] n1828;
wire     [31:0] n1829;
wire     [31:0] n1830;
wire     [31:0] n1831;
wire     [31:0] n1832;
wire     [31:0] n1833;
wire     [31:0] n1834;
wire     [31:0] n1835;
wire     [31:0] n1836;
wire     [31:0] n1837;
wire     [31:0] n1838;
wire     [31:0] n1839;
wire     [31:0] n1840;
wire     [31:0] n1841;
wire     [31:0] n1842;
wire     [31:0] n1843;
wire     [31:0] n1844;
wire     [31:0] n1845;
wire     [31:0] n1846;
wire     [31:0] n1847;
wire     [31:0] n1848;
wire     [31:0] n1849;
wire     [31:0] n1850;
wire     [31:0] n1851;
wire     [31:0] n1852;
wire     [31:0] n1853;
wire     [31:0] n1854;
wire     [31:0] n1855;
wire     [31:0] n1856;
wire     [31:0] n1857;
wire     [31:0] n1858;
wire     [31:0] n1859;
wire     [31:0] n1860;
wire            n1861;
wire     [31:0] n1862;
wire     [31:0] n1863;
wire     [31:0] n1864;
wire     [31:0] n1865;
wire     [31:0] n1866;
wire     [31:0] n1867;
wire     [31:0] n1868;
wire     [31:0] n1869;
wire     [31:0] n1870;
wire     [31:0] n1871;
wire     [31:0] n1872;
wire     [31:0] n1873;
wire     [31:0] n1874;
wire     [31:0] n1875;
wire     [31:0] n1876;
wire     [31:0] n1877;
wire     [31:0] n1878;
wire     [31:0] n1879;
wire     [31:0] n1880;
wire     [31:0] n1881;
wire     [31:0] n1882;
wire     [31:0] n1883;
wire     [31:0] n1884;
wire     [31:0] n1885;
wire     [31:0] n1886;
wire     [31:0] n1887;
wire     [31:0] n1888;
wire     [31:0] n1889;
wire     [31:0] n1890;
wire     [31:0] n1891;
wire     [31:0] n1892;
wire     [31:0] n1893;
wire     [31:0] n1894;
wire     [31:0] n1895;
wire     [31:0] n1896;
wire     [31:0] n1897;
wire     [31:0] n1898;
wire     [31:0] n1899;
wire     [31:0] n1900;
wire     [31:0] n1901;
wire     [31:0] n1902;
wire     [31:0] n1903;
wire     [31:0] n1904;
wire     [31:0] n1905;
wire     [31:0] n1906;
wire     [31:0] n1907;
wire     [31:0] n1908;
wire     [31:0] n1909;
wire     [31:0] n1910;
wire     [31:0] n1911;
wire     [31:0] n1912;
wire     [31:0] n1913;
wire     [31:0] n1914;
wire     [31:0] n1915;
wire     [31:0] n1916;
wire            n1917;
wire     [31:0] n1918;
wire     [31:0] n1919;
wire     [31:0] n1920;
wire     [31:0] n1921;
wire     [31:0] n1922;
wire     [31:0] n1923;
wire     [31:0] n1924;
wire     [31:0] n1925;
wire     [31:0] n1926;
wire     [31:0] n1927;
wire     [31:0] n1928;
wire     [31:0] n1929;
wire     [31:0] n1930;
wire     [31:0] n1931;
wire     [31:0] n1932;
wire     [31:0] n1933;
wire     [31:0] n1934;
wire     [31:0] n1935;
wire     [31:0] n1936;
wire     [31:0] n1937;
wire     [31:0] n1938;
wire     [31:0] n1939;
wire     [31:0] n1940;
wire     [31:0] n1941;
wire     [31:0] n1942;
wire     [31:0] n1943;
wire     [31:0] n1944;
wire     [31:0] n1945;
wire     [31:0] n1946;
wire     [31:0] n1947;
wire     [31:0] n1948;
wire     [31:0] n1949;
wire     [31:0] n1950;
wire     [31:0] n1951;
wire     [31:0] n1952;
wire     [31:0] n1953;
wire     [31:0] n1954;
wire     [31:0] n1955;
wire     [31:0] n1956;
wire     [31:0] n1957;
wire     [31:0] n1958;
wire     [31:0] n1959;
wire     [31:0] n1960;
wire     [31:0] n1961;
wire     [31:0] n1962;
wire     [31:0] n1963;
wire     [31:0] n1964;
wire     [31:0] n1965;
wire     [31:0] n1966;
wire     [31:0] n1967;
wire     [31:0] n1968;
wire     [31:0] n1969;
wire     [31:0] n1970;
wire     [31:0] n1971;
wire            n1972;
wire     [31:0] n1973;
wire     [31:0] n1974;
wire     [31:0] n1975;
wire     [31:0] n1976;
wire     [31:0] n1977;
wire     [31:0] n1978;
wire     [31:0] n1979;
wire     [31:0] n1980;
wire     [31:0] n1981;
wire     [31:0] n1982;
wire     [31:0] n1983;
wire     [31:0] n1984;
wire     [31:0] n1985;
wire     [31:0] n1986;
wire     [31:0] n1987;
wire     [31:0] n1988;
wire     [31:0] n1989;
wire     [31:0] n1990;
wire     [31:0] n1991;
wire     [31:0] n1992;
wire     [31:0] n1993;
wire     [31:0] n1994;
wire     [31:0] n1995;
wire     [31:0] n1996;
wire     [31:0] n1997;
wire     [31:0] n1998;
wire     [31:0] n1999;
wire     [31:0] n2000;
wire     [31:0] n2001;
wire     [31:0] n2002;
wire     [31:0] n2003;
wire     [31:0] n2004;
wire     [31:0] n2005;
wire     [31:0] n2006;
wire     [31:0] n2007;
wire     [31:0] n2008;
wire     [31:0] n2009;
wire     [31:0] n2010;
wire     [31:0] n2011;
wire     [31:0] n2012;
wire     [31:0] n2013;
wire     [31:0] n2014;
wire     [31:0] n2015;
wire     [31:0] n2016;
wire     [31:0] n2017;
wire     [31:0] n2018;
wire     [31:0] n2019;
wire     [31:0] n2020;
wire     [31:0] n2021;
wire     [31:0] n2022;
wire     [31:0] n2023;
wire     [31:0] n2024;
wire     [31:0] n2025;
wire     [31:0] n2026;
wire            n2027;
wire     [31:0] n2028;
wire     [31:0] n2029;
wire     [31:0] n2030;
wire     [31:0] n2031;
wire     [31:0] n2032;
wire     [31:0] n2033;
wire     [31:0] n2034;
wire     [31:0] n2035;
wire     [31:0] n2036;
wire     [31:0] n2037;
wire     [31:0] n2038;
wire     [31:0] n2039;
wire     [31:0] n2040;
wire     [31:0] n2041;
wire     [31:0] n2042;
wire     [31:0] n2043;
wire     [31:0] n2044;
wire     [31:0] n2045;
wire     [31:0] n2046;
wire     [31:0] n2047;
wire     [31:0] n2048;
wire     [31:0] n2049;
wire     [31:0] n2050;
wire     [31:0] n2051;
wire     [31:0] n2052;
wire     [31:0] n2053;
wire     [31:0] n2054;
wire     [31:0] n2055;
wire     [31:0] n2056;
wire     [31:0] n2057;
wire     [31:0] n2058;
wire     [31:0] n2059;
wire     [31:0] n2060;
wire     [31:0] n2061;
wire     [31:0] n2062;
wire     [31:0] n2063;
wire     [31:0] n2064;
wire     [31:0] n2065;
wire     [31:0] n2066;
wire     [31:0] n2067;
wire     [31:0] n2068;
wire     [31:0] n2069;
wire     [31:0] n2070;
wire     [31:0] n2071;
wire     [31:0] n2072;
wire     [31:0] n2073;
wire     [31:0] n2074;
wire     [31:0] n2075;
wire     [31:0] n2076;
wire     [31:0] n2077;
wire     [31:0] n2078;
wire     [31:0] n2079;
wire     [31:0] n2080;
wire     [31:0] n2081;
wire     [31:0] mem_addr0;
wire     [31:0] mem_data0;
wire            n2082;
wire            n2083;
wire            n2084;
wire            n2085;
wire            n2086;
wire            n2087;
wire     [11:0] n2088;
wire     [31:0] n2089;
wire     [31:0] n2090;
wire     [29:0] n2091;
wire     [31:0] n2092;
wire     [31:0] n2093;
wire      [1:0] n2094;
wire     [31:0] n2095;
wire     [31:0] n2096;
wire     [31:0] n2097;
wire     [31:0] n2098;
wire     [31:0] n2099;
wire     [31:0] n2100;
wire     [31:0] n2101;
wire     [31:0] n2102;
wire            n2103;
wire     [31:0] n2104;
wire     [31:0] n2105;
wire     [31:0] n2106;
wire     [31:0] n2107;
wire     [31:0] n2108;
wire     [31:0] n2109;
wire     [31:0] n2110;
wire     [31:0] n2111;
wire     [31:0] n2112;
wire     [31:0] n2113;
wire     [31:0] n2114;
wire     [31:0] n2115;
//reg     [31:0] mem;
wire clk;
wire rst;
wire step;
assign n0 = pc[31:2] ;
assign n1 =  {2'd0 , n0}  ;
//assign n2 =  (  mem [ n1 ] )  ;
assign mem_raddr0 = n1;
assign n2 = mem_rdata0;

assign n3 = n2[6:0] ;
assign n4 =  ( n3 ) == ( 7'd103 )  ;
assign n5 = n2[14:12] ;
assign n6 =  ( n5 ) == ( 3'd0 )  ;
assign n7 =  ( n4 ) & ( n6 )  ;
assign n8 = n2[19:15] ;
assign n9 =  ( n8 ) == ( 5'd31 )  ;
assign n10 =  ( n8 ) == ( 5'd30 )  ;
assign n11 =  ( n8 ) == ( 5'd29 )  ;
assign n12 =  ( n8 ) == ( 5'd28 )  ;
assign n13 =  ( n8 ) == ( 5'd27 )  ;
assign n14 =  ( n8 ) == ( 5'd26 )  ;
assign n15 =  ( n8 ) == ( 5'd25 )  ;
assign n16 =  ( n8 ) == ( 5'd24 )  ;
assign n17 =  ( n8 ) == ( 5'd23 )  ;
assign n18 =  ( n8 ) == ( 5'd22 )  ;
assign n19 =  ( n8 ) == ( 5'd21 )  ;
assign n20 =  ( n8 ) == ( 5'd20 )  ;
assign n21 =  ( n8 ) == ( 5'd19 )  ;
assign n22 =  ( n8 ) == ( 5'd18 )  ;
assign n23 =  ( n8 ) == ( 5'd17 )  ;
assign n24 =  ( n8 ) == ( 5'd16 )  ;
assign n25 =  ( n8 ) == ( 5'd15 )  ;
assign n26 =  ( n8 ) == ( 5'd14 )  ;
assign n27 =  ( n8 ) == ( 5'd13 )  ;
assign n28 =  ( n8 ) == ( 5'd12 )  ;
assign n29 =  ( n8 ) == ( 5'd11 )  ;
assign n30 =  ( n8 ) == ( 5'd10 )  ;
assign n31 =  ( n8 ) == ( 5'd9 )  ;
assign n32 =  ( n8 ) == ( 5'd8 )  ;
assign n33 =  ( n8 ) == ( 5'd7 )  ;
assign n34 =  ( n8 ) == ( 5'd6 )  ;
assign n35 =  ( n8 ) == ( 5'd5 )  ;
assign n36 =  ( n8 ) == ( 5'd4 )  ;
assign n37 =  ( n8 ) == ( 5'd3 )  ;
assign n38 =  ( n8 ) == ( 5'd2 )  ;
assign n39 =  ( n8 ) == ( 5'd1 )  ;
assign n40 =  ( n39 ) ? ( x1 ) : ( x0 ) ;
assign n41 =  ( n38 ) ? ( x2 ) : ( n40 ) ;
assign n42 =  ( n37 ) ? ( x3 ) : ( n41 ) ;
assign n43 =  ( n36 ) ? ( x4 ) : ( n42 ) ;
assign n44 =  ( n35 ) ? ( x5 ) : ( n43 ) ;
assign n45 =  ( n34 ) ? ( x6 ) : ( n44 ) ;
assign n46 =  ( n33 ) ? ( x7 ) : ( n45 ) ;
assign n47 =  ( n32 ) ? ( x8 ) : ( n46 ) ;
assign n48 =  ( n31 ) ? ( x9 ) : ( n47 ) ;
assign n49 =  ( n30 ) ? ( x10 ) : ( n48 ) ;
assign n50 =  ( n29 ) ? ( x11 ) : ( n49 ) ;
assign n51 =  ( n28 ) ? ( x12 ) : ( n50 ) ;
assign n52 =  ( n27 ) ? ( x13 ) : ( n51 ) ;
assign n53 =  ( n26 ) ? ( x14 ) : ( n52 ) ;
assign n54 =  ( n25 ) ? ( x15 ) : ( n53 ) ;
assign n55 =  ( n24 ) ? ( x16 ) : ( n54 ) ;
assign n56 =  ( n23 ) ? ( x17 ) : ( n55 ) ;
assign n57 =  ( n22 ) ? ( x18 ) : ( n56 ) ;
assign n58 =  ( n21 ) ? ( x19 ) : ( n57 ) ;
assign n59 =  ( n20 ) ? ( x20 ) : ( n58 ) ;
assign n60 =  ( n19 ) ? ( x21 ) : ( n59 ) ;
assign n61 =  ( n18 ) ? ( x22 ) : ( n60 ) ;
assign n62 =  ( n17 ) ? ( x23 ) : ( n61 ) ;
assign n63 =  ( n16 ) ? ( x24 ) : ( n62 ) ;
assign n64 =  ( n15 ) ? ( x25 ) : ( n63 ) ;
assign n65 =  ( n14 ) ? ( x26 ) : ( n64 ) ;
assign n66 =  ( n13 ) ? ( x27 ) : ( n65 ) ;
assign n67 =  ( n12 ) ? ( x28 ) : ( n66 ) ;
assign n68 =  ( n11 ) ? ( x29 ) : ( n67 ) ;
assign n69 =  ( n10 ) ? ( x30 ) : ( n68 ) ;
assign n70 =  ( n9 ) ? ( x31 ) : ( n69 ) ;
assign n71 = n2[31:20] ;
assign n72 =  { {20{n71[11] }  }, n71}  ;
assign n73 =  ( n70 ) + ( n72 )  ;
assign n74 =  ( n73 ) & ( 32'd4294967294 )  ;
assign n75 =  ( n3 ) == ( 7'd111 )  ;
assign n76 = n2[31:31] ;
assign n77 = n2[19:12] ;
assign n78 = n2[20:20] ;
assign n79 = n2[30:21] ;
assign n80 =  { ( n79 ) , ( 1'd0 ) }  ;
assign n81 =  { ( n78 ) , ( n80 ) }  ;
assign n82 =  { ( n77 ) , ( n81 ) }  ;
assign n83 =  { ( n76 ) , ( n82 ) }  ;
assign n84 =  { {11{n83[20] }  }, n83}  ;
assign n85 =  ( pc ) + ( n84 )  ;
assign n86 =  ( n3 ) == ( 7'd99 )  ;
assign n87 =  ( n5 ) == ( 3'd7 )  ;
assign n88 =  ( n86 ) & ( n87 )  ;
assign n89 = n2[24:20] ;
assign n90 =  ( n89 ) == ( 5'd31 )  ;
assign n91 =  ( n89 ) == ( 5'd30 )  ;
assign n92 =  ( n89 ) == ( 5'd29 )  ;
assign n93 =  ( n89 ) == ( 5'd28 )  ;
assign n94 =  ( n89 ) == ( 5'd27 )  ;
assign n95 =  ( n89 ) == ( 5'd26 )  ;
assign n96 =  ( n89 ) == ( 5'd25 )  ;
assign n97 =  ( n89 ) == ( 5'd24 )  ;
assign n98 =  ( n89 ) == ( 5'd23 )  ;
assign n99 =  ( n89 ) == ( 5'd22 )  ;
assign n100 =  ( n89 ) == ( 5'd21 )  ;
assign n101 =  ( n89 ) == ( 5'd20 )  ;
assign n102 =  ( n89 ) == ( 5'd19 )  ;
assign n103 =  ( n89 ) == ( 5'd18 )  ;
assign n104 =  ( n89 ) == ( 5'd17 )  ;
assign n105 =  ( n89 ) == ( 5'd16 )  ;
assign n106 =  ( n89 ) == ( 5'd15 )  ;
assign n107 =  ( n89 ) == ( 5'd14 )  ;
assign n108 =  ( n89 ) == ( 5'd13 )  ;
assign n109 =  ( n89 ) == ( 5'd12 )  ;
assign n110 =  ( n89 ) == ( 5'd11 )  ;
assign n111 =  ( n89 ) == ( 5'd10 )  ;
assign n112 =  ( n89 ) == ( 5'd9 )  ;
assign n113 =  ( n89 ) == ( 5'd8 )  ;
assign n114 =  ( n89 ) == ( 5'd7 )  ;
assign n115 =  ( n89 ) == ( 5'd6 )  ;
assign n116 =  ( n89 ) == ( 5'd5 )  ;
assign n117 =  ( n89 ) == ( 5'd4 )  ;
assign n118 =  ( n89 ) == ( 5'd3 )  ;
assign n119 =  ( n89 ) == ( 5'd2 )  ;
assign n120 =  ( n89 ) == ( 5'd1 )  ;
assign n121 =  ( n120 ) ? ( x1 ) : ( x0 ) ;
assign n122 =  ( n119 ) ? ( x2 ) : ( n121 ) ;
assign n123 =  ( n118 ) ? ( x3 ) : ( n122 ) ;
assign n124 =  ( n117 ) ? ( x4 ) : ( n123 ) ;
assign n125 =  ( n116 ) ? ( x5 ) : ( n124 ) ;
assign n126 =  ( n115 ) ? ( x6 ) : ( n125 ) ;
assign n127 =  ( n114 ) ? ( x7 ) : ( n126 ) ;
assign n128 =  ( n113 ) ? ( x8 ) : ( n127 ) ;
assign n129 =  ( n112 ) ? ( x9 ) : ( n128 ) ;
assign n130 =  ( n111 ) ? ( x10 ) : ( n129 ) ;
assign n131 =  ( n110 ) ? ( x11 ) : ( n130 ) ;
assign n132 =  ( n109 ) ? ( x12 ) : ( n131 ) ;
assign n133 =  ( n108 ) ? ( x13 ) : ( n132 ) ;
assign n134 =  ( n107 ) ? ( x14 ) : ( n133 ) ;
assign n135 =  ( n106 ) ? ( x15 ) : ( n134 ) ;
assign n136 =  ( n105 ) ? ( x16 ) : ( n135 ) ;
assign n137 =  ( n104 ) ? ( x17 ) : ( n136 ) ;
assign n138 =  ( n103 ) ? ( x18 ) : ( n137 ) ;
assign n139 =  ( n102 ) ? ( x19 ) : ( n138 ) ;
assign n140 =  ( n101 ) ? ( x20 ) : ( n139 ) ;
assign n141 =  ( n100 ) ? ( x21 ) : ( n140 ) ;
assign n142 =  ( n99 ) ? ( x22 ) : ( n141 ) ;
assign n143 =  ( n98 ) ? ( x23 ) : ( n142 ) ;
assign n144 =  ( n97 ) ? ( x24 ) : ( n143 ) ;
assign n145 =  ( n96 ) ? ( x25 ) : ( n144 ) ;
assign n146 =  ( n95 ) ? ( x26 ) : ( n145 ) ;
assign n147 =  ( n94 ) ? ( x27 ) : ( n146 ) ;
assign n148 =  ( n93 ) ? ( x28 ) : ( n147 ) ;
assign n149 =  ( n92 ) ? ( x29 ) : ( n148 ) ;
assign n150 =  ( n91 ) ? ( x30 ) : ( n149 ) ;
assign n151 =  ( n90 ) ? ( x31 ) : ( n150 ) ;
assign n152 =  ( n70 ) >= ( n151 )  ;
assign n153 = n2[7:7] ;
assign n154 = n2[30:25] ;
assign n155 = n2[11:8] ;
assign n156 =  { ( n155 ) , ( 1'd0 ) }  ;
assign n157 =  { ( n154 ) , ( n156 ) }  ;
assign n158 =  { ( n153 ) , ( n157 ) }  ;
assign n159 =  { ( n76 ) , ( n158 ) }  ;
assign n160 =  { {19{n159[12] }  }, n159}  ;
assign n161 =  ( pc ) + ( n160 )  ;
assign n162 =  ( pc ) + ( 32'd4 )  ;
assign n163 =  ( n152 ) ? ( n161 ) : ( n162 ) ;
assign n164 =  ( n5 ) == ( 3'd5 )  ;
assign n165 =  ( n86 ) & ( n164 )  ;
assign n166 =  $signed( n70 ) >= $signed( n151 )  ;
assign n167 =  ( n166 ) ? ( n161 ) : ( n162 ) ;
assign n168 =  ( n5 ) == ( 3'd6 )  ;
assign n169 =  ( n86 ) & ( n168 )  ;
assign n170 =  ( n70 ) < ( n151 )  ;
assign n171 =  ( n170 ) ? ( n161 ) : ( n162 ) ;
assign n172 =  ( n5 ) == ( 3'd4 )  ;
assign n173 =  ( n86 ) & ( n172 )  ;
assign n174 =  $signed( n70 ) < $signed( n151 )  ;
assign n175 =  ( n174 ) ? ( n161 ) : ( n162 ) ;
assign n176 =  ( n5 ) == ( 3'd1 )  ;
assign n177 =  ( n86 ) & ( n176 )  ;
assign n178 =  ( n70 ) != ( n151 )  ;
assign n179 =  ( n178 ) ? ( n161 ) : ( n162 ) ;
assign n180 =  ( n86 ) & ( n6 )  ;
assign n181 =  ( n70 ) == ( n151 )  ;
assign n182 =  ( n181 ) ? ( n161 ) : ( n162 ) ;
assign n183 =  ( n3 ) == ( 7'd51 )  ;
assign n184 =  ( n183 ) & ( n164 )  ;
assign n185 = n2[31:25] ;
assign n186 =  ( n185 ) == ( 7'd32 )  ;
assign n187 =  ( n184 ) & ( n186 )  ;
assign n188 =  ( n183 ) & ( n6 )  ;
assign n189 =  ( n188 ) & ( n186 )  ;
assign n190 =  ( n185 ) == ( 7'd0 )  ;
assign n191 =  ( n184 ) & ( n190 )  ;
assign n192 =  ( n183 ) & ( n176 )  ;
assign n193 =  ( n192 ) & ( n190 )  ;
assign n194 =  ( n183 ) & ( n172 )  ;
assign n195 =  ( n194 ) & ( n190 )  ;
assign n196 =  ( n183 ) & ( n168 )  ;
assign n197 =  ( n196 ) & ( n190 )  ;
assign n198 =  ( n183 ) & ( n87 )  ;
assign n199 =  ( n198 ) & ( n190 )  ;
assign n200 =  ( n5 ) == ( 3'd3 )  ;
assign n201 =  ( n183 ) & ( n200 )  ;
assign n202 =  ( n201 ) & ( n190 )  ;
assign n203 =  ( n5 ) == ( 3'd2 )  ;
assign n204 =  ( n183 ) & ( n203 )  ;
assign n205 =  ( n204 ) & ( n190 )  ;
assign n206 =  ( n188 ) & ( n190 )  ;
assign n207 =  ( n3 ) == ( 7'd19 )  ;
assign n208 =  ( n207 ) & ( n164 )  ;
assign n209 =  ( n208 ) & ( n186 )  ;
assign n210 =  ( n208 ) & ( n190 )  ;
assign n211 =  ( n207 ) & ( n176 )  ;
assign n212 =  ( n211 ) & ( n190 )  ;
assign n213 =  ( n207 ) & ( n172 )  ;
assign n214 =  ( n207 ) & ( n168 )  ;
assign n215 =  ( n207 ) & ( n87 )  ;
assign n216 =  ( n207 ) & ( n200 )  ;
assign n217 =  ( n207 ) & ( n203 )  ;
assign n218 =  ( n207 ) & ( n6 )  ;
assign n219 =  ( n3 ) == ( 7'd23 )  ;
assign n220 =  ( n3 ) == ( 7'd55 )  ;
assign n221 =  ( n3 ) == ( 7'd35 )  ;
assign n222 =  ( n221 ) & ( n203 )  ;
assign n223 =  ( n221 ) & ( n176 )  ;
assign n224 =  ( n221 ) & ( n6 )  ;
assign n225 =  ( n3 ) == ( 7'd3 )  ;
assign n226 =  ( n225 ) & ( n164 )  ;
assign n227 =  ( n225 ) & ( n172 )  ;
assign n228 =  ( n225 ) & ( n6 )  ;
assign n229 =  ( n225 ) & ( n176 )  ;
assign n230 =  ( n225 ) & ( n203 )  ;
assign n231 =  ( n229 ) | ( n230 )  ;
assign n232 =  ( n228 ) | ( n231 )  ;
assign n233 =  ( n227 ) | ( n232 )  ;
assign n234 =  ( n226 ) | ( n233 )  ;
assign n235 =  ( n224 ) | ( n234 )  ;
assign n236 =  ( n223 ) | ( n235 )  ;
assign n237 =  ( n222 ) | ( n236 )  ;
assign n238 =  ( n220 ) | ( n237 )  ;
assign n239 =  ( n219 ) | ( n238 )  ;
assign n240 =  ( n218 ) | ( n239 )  ;
assign n241 =  ( n217 ) | ( n240 )  ;
assign n242 =  ( n216 ) | ( n241 )  ;
assign n243 =  ( n215 ) | ( n242 )  ;
assign n244 =  ( n214 ) | ( n243 )  ;
assign n245 =  ( n213 ) | ( n244 )  ;
assign n246 =  ( n212 ) | ( n245 )  ;
assign n247 =  ( n210 ) | ( n246 )  ;
assign n248 =  ( n209 ) | ( n247 )  ;
assign n249 =  ( n206 ) | ( n248 )  ;
assign n250 =  ( n205 ) | ( n249 )  ;
assign n251 =  ( n202 ) | ( n250 )  ;
assign n252 =  ( n199 ) | ( n251 )  ;
assign n253 =  ( n197 ) | ( n252 )  ;
assign n254 =  ( n195 ) | ( n253 )  ;
assign n255 =  ( n193 ) | ( n254 )  ;
assign n256 =  ( n191 ) | ( n255 )  ;
assign n257 =  ( n189 ) | ( n256 )  ;
assign n258 =  ( n187 ) | ( n257 )  ;
assign n259 =  ( n258 ) ? ( n162 ) : ( pc ) ;
assign n260 =  ( n180 ) ? ( n182 ) : ( n259 ) ;
assign n261 =  ( n177 ) ? ( n179 ) : ( n260 ) ;
assign n262 =  ( n173 ) ? ( n175 ) : ( n261 ) ;
assign n263 =  ( n169 ) ? ( n171 ) : ( n262 ) ;
assign n264 =  ( n165 ) ? ( n167 ) : ( n263 ) ;
assign n265 =  ( n88 ) ? ( n163 ) : ( n264 ) ;
assign n266 =  ( n75 ) ? ( n85 ) : ( n265 ) ;
assign n267 =  ( n7 ) ? ( n74 ) : ( n266 ) ;
assign n268 =  ( n180 ) | ( n239 )  ;
assign n269 =  ( n177 ) | ( n268 )  ;
assign n270 =  ( n173 ) | ( n269 )  ;
assign n271 =  ( n169 ) | ( n270 )  ;
assign n272 =  ( n165 ) | ( n271 )  ;
assign n273 =  ( n88 ) | ( n272 )  ;
assign n274 =  ( n75 ) | ( n273 )  ;
assign n275 =  ( n7 ) | ( n274 )  ;
assign n276 =  ( n218 ) | ( n275 )  ;
assign n277 =  ( n217 ) | ( n276 )  ;
assign n278 =  ( n216 ) | ( n277 )  ;
assign n279 =  ( n215 ) | ( n278 )  ;
assign n280 =  ( n214 ) | ( n279 )  ;
assign n281 =  ( n213 ) | ( n280 )  ;
assign n282 =  ( n212 ) | ( n281 )  ;
assign n283 =  ( n210 ) | ( n282 )  ;
assign n284 =  ( n209 ) | ( n283 )  ;
assign n285 =  ( n206 ) | ( n284 )  ;
assign n286 =  ( n205 ) | ( n285 )  ;
assign n287 =  ( n202 ) | ( n286 )  ;
assign n288 =  ( n199 ) | ( n287 )  ;
assign n289 =  ( n197 ) | ( n288 )  ;
assign n290 =  ( n195 ) | ( n289 )  ;
assign n291 =  ( n193 ) | ( n290 )  ;
assign n292 =  ( n191 ) | ( n291 )  ;
assign n293 =  ( n189 ) | ( n292 )  ;
assign n294 =  ( n187 ) | ( n293 )  ;
assign n295 =  ( n294 ) ? ( 32'd0 ) : ( x0 ) ;
assign n296 = n2[11:7] ;
assign n297 =  ( n296 ) == ( 5'd1 )  ;
assign n298 = n151[4:0] ;
assign n299 =  {27'd0 , n298}  ;
assign n300 =  ( $signed( n70 ) >>> ( n299 ))  ;
assign n301 =  ( n297 ) ? ( n300 ) : ( x1 ) ;
assign n302 =  ( n70 ) - ( n151 )  ;
assign n303 =  ( n297 ) ? ( n302 ) : ( x1 ) ;
assign n304 =  ( ( n70 ) >> ( n299 ))  ;
assign n305 =  ( n297 ) ? ( n304 ) : ( x1 ) ;
assign n306 =  ( n70 ) << ( n299 )  ;
assign n307 =  ( n297 ) ? ( n306 ) : ( x1 ) ;
assign n308 =  ( n70 ) ^ ( n151 )  ;
assign n309 =  ( n297 ) ? ( n308 ) : ( x1 ) ;
assign n310 =  ( n70 ) | ( n151 )  ;
assign n311 =  ( n297 ) ? ( n310 ) : ( x1 ) ;
assign n312 =  ( n70 ) & ( n151 )  ;
assign n313 =  ( n297 ) ? ( n312 ) : ( x1 ) ;
assign n314 =  ( n170 ) ? ( 32'd1 ) : ( 32'd0 ) ;
assign n315 =  ( n297 ) ? ( n314 ) : ( x1 ) ;
assign n316 =  ( n174 ) ? ( 32'd1 ) : ( 32'd0 ) ;
assign n317 =  ( n297 ) ? ( n316 ) : ( x1 ) ;
assign n318 =  ( n70 ) + ( n151 )  ;
assign n319 =  ( n297 ) ? ( n318 ) : ( x1 ) ;
assign n320 =  {27'd0 , n89}  ;
assign n321 =  ( $signed( n70 ) >>> ( n320 ))  ;
assign n322 =  ( n297 ) ? ( n321 ) : ( x1 ) ;
assign n323 =  ( ( n70 ) >> ( n320 ))  ;
assign n324 =  ( n297 ) ? ( n323 ) : ( x1 ) ;
assign n325 =  ( n70 ) << ( n320 )  ;
assign n326 =  ( n297 ) ? ( n325 ) : ( x1 ) ;
assign n327 = n72 ;
assign n328 =  ( n70 ) ^ ( n327 )  ;
assign n329 =  ( n297 ) ? ( n328 ) : ( x1 ) ;
assign n330 = n72 ;
assign n331 =  ( n70 ) | ( n330 )  ;
assign n332 =  ( n297 ) ? ( n331 ) : ( x1 ) ;
assign n333 =  ( n70 ) & ( n327 )  ;
assign n334 =  ( n297 ) ? ( n333 ) : ( x1 ) ;
assign n335 =  ( n70 ) < ( n330 )  ;
assign n336 =  ( n335 ) ? ( 32'd1 ) : ( 32'd0 ) ;
assign n337 =  ( n297 ) ? ( n336 ) : ( x1 ) ;
assign n338 =  $signed( n70 ) < $signed( n327 )  ;
assign n339 =  ( n338 ) ? ( 32'd1 ) : ( 32'd0 ) ;
assign n340 =  ( n297 ) ? ( n339 ) : ( x1 ) ;
assign n341 =  ( n70 ) + ( n327 )  ;
assign n342 =  ( n297 ) ? ( n341 ) : ( x1 ) ;
assign n343 =  ( n7 ) | ( n75 )  ;
assign n344 =  ( n297 ) ? ( n162 ) : ( x1 ) ;
assign n345 = n2[31:12] ;
assign n346 =  { ( n345 ) , ( 12'd0 ) }  ;
assign n347 =  ( n346 ) + ( pc )  ;
assign n348 =  ( n297 ) ? ( n347 ) : ( x1 ) ;
assign n349 =  ( n297 ) ? ( n346 ) : ( x1 ) ;
assign n350 = n73[1:0] ;
assign n351 =  ( n350 ) == ( 2'd0 )  ;
assign n352 = n73[31:2] ;
assign n353 =  {2'd0 , n352}  ;
//assign n354 =  (  mem [ n353 ] )  ;
assign mem_raddr1 = n353;
assign n354 = mem_rdata1;

assign n355 = n354[15:0] ;
assign n356 =  {16'd0 , n355}  ;
assign n357 =  ( n350 ) == ( 2'd1 )  ;
assign n358 = n354[15:8] ;
assign n359 =  {24'd0 , n358}  ;
assign n360 =  ( n350 ) == ( 2'd2 )  ;
assign n361 = n354[31:16] ;
assign n362 =  {16'd0 , n361}  ;
assign n363 =  ( n350 ) == ( 2'd3 )  ;
assign n364 = n354[31:24] ;
assign n365 =  {24'd0 , n364}  ;
assign n366 = n354[31:0] ;
assign n367 =  ( n363 ) ? ( n365 ) : ( n366 ) ;
assign n368 =  ( n360 ) ? ( n362 ) : ( n367 ) ;
assign n369 =  ( n357 ) ? ( n359 ) : ( n368 ) ;
assign n370 =  ( n351 ) ? ( n356 ) : ( n369 ) ;
assign n371 =  ( n297 ) ? ( n370 ) : ( x1 ) ;
assign n372 = n354[7:0] ;
assign n373 =  {24'd0 , n372}  ;
assign n374 = n354[23:16] ;
assign n375 =  {24'd0 , n374}  ;
assign n376 =  ( n360 ) ? ( n375 ) : ( n367 ) ;
assign n377 =  ( n357 ) ? ( n359 ) : ( n376 ) ;
assign n378 =  ( n351 ) ? ( n373 ) : ( n377 ) ;
assign n379 =  ( n297 ) ? ( n378 ) : ( x1 ) ;
assign n380 =  { {24{n372[7] }  }, n372}  ;
assign n381 =  { {24{n358[7] }  }, n358}  ;
assign n382 =  { {24{n374[7] }  }, n374}  ;
assign n383 =  { {24{n364[7] }  }, n364}  ;
assign n384 =  ( n363 ) ? ( n383 ) : ( n366 ) ;
assign n385 =  ( n360 ) ? ( n382 ) : ( n384 ) ;
assign n386 =  ( n357 ) ? ( n381 ) : ( n385 ) ;
assign n387 =  ( n351 ) ? ( n380 ) : ( n386 ) ;
assign n388 =  ( n297 ) ? ( n387 ) : ( x1 ) ;
assign n389 =  { {16{n355[15] }  }, n355}  ;
assign n390 =  { {16{n361[15] }  }, n361}  ;
assign n391 =  ( n360 ) ? ( n390 ) : ( n367 ) ;
assign n392 =  ( n357 ) ? ( n359 ) : ( n391 ) ;
assign n393 =  ( n351 ) ? ( n389 ) : ( n392 ) ;
assign n394 =  ( n297 ) ? ( n393 ) : ( x1 ) ;
assign n395 =  ( n351 ) ? ( n366 ) : ( n377 ) ;
assign n396 =  ( n297 ) ? ( n395 ) : ( x1 ) ;
assign n397 =  ( n230 ) ? ( n396 ) : ( x1 ) ;
assign n398 =  ( n229 ) ? ( n394 ) : ( n397 ) ;
assign n399 =  ( n228 ) ? ( n388 ) : ( n398 ) ;
assign n400 =  ( n227 ) ? ( n379 ) : ( n399 ) ;
assign n401 =  ( n226 ) ? ( n371 ) : ( n400 ) ;
assign n402 =  ( n220 ) ? ( n349 ) : ( n401 ) ;
assign n403 =  ( n219 ) ? ( n348 ) : ( n402 ) ;
assign n404 =  ( n343 ) ? ( n344 ) : ( n403 ) ;
assign n405 =  ( n218 ) ? ( n342 ) : ( n404 ) ;
assign n406 =  ( n217 ) ? ( n340 ) : ( n405 ) ;
assign n407 =  ( n216 ) ? ( n337 ) : ( n406 ) ;
assign n408 =  ( n215 ) ? ( n334 ) : ( n407 ) ;
assign n409 =  ( n214 ) ? ( n332 ) : ( n408 ) ;
assign n410 =  ( n213 ) ? ( n329 ) : ( n409 ) ;
assign n411 =  ( n212 ) ? ( n326 ) : ( n410 ) ;
assign n412 =  ( n210 ) ? ( n324 ) : ( n411 ) ;
assign n413 =  ( n209 ) ? ( n322 ) : ( n412 ) ;
assign n414 =  ( n206 ) ? ( n319 ) : ( n413 ) ;
assign n415 =  ( n205 ) ? ( n317 ) : ( n414 ) ;
assign n416 =  ( n202 ) ? ( n315 ) : ( n415 ) ;
assign n417 =  ( n199 ) ? ( n313 ) : ( n416 ) ;
assign n418 =  ( n197 ) ? ( n311 ) : ( n417 ) ;
assign n419 =  ( n195 ) ? ( n309 ) : ( n418 ) ;
assign n420 =  ( n193 ) ? ( n307 ) : ( n419 ) ;
assign n421 =  ( n191 ) ? ( n305 ) : ( n420 ) ;
assign n422 =  ( n189 ) ? ( n303 ) : ( n421 ) ;
assign n423 =  ( n187 ) ? ( n301 ) : ( n422 ) ;
assign n424 =  ( n296 ) == ( 5'd10 )  ;
assign n425 =  ( n424 ) ? ( n300 ) : ( x10 ) ;
assign n426 =  ( n424 ) ? ( n302 ) : ( x10 ) ;
assign n427 =  ( n424 ) ? ( n304 ) : ( x10 ) ;
assign n428 =  ( n424 ) ? ( n306 ) : ( x10 ) ;
assign n429 =  ( n424 ) ? ( n308 ) : ( x10 ) ;
assign n430 =  ( n424 ) ? ( n310 ) : ( x10 ) ;
assign n431 =  ( n424 ) ? ( n312 ) : ( x10 ) ;
assign n432 =  ( n424 ) ? ( n314 ) : ( x10 ) ;
assign n433 =  ( n424 ) ? ( n316 ) : ( x10 ) ;
assign n434 =  ( n424 ) ? ( n318 ) : ( x10 ) ;
assign n435 =  ( n424 ) ? ( n321 ) : ( x10 ) ;
assign n436 =  ( n424 ) ? ( n323 ) : ( x10 ) ;
assign n437 =  ( n424 ) ? ( n325 ) : ( x10 ) ;
assign n438 =  ( n424 ) ? ( n328 ) : ( x10 ) ;
assign n439 =  ( n70 ) | ( n327 )  ;
assign n440 =  ( n424 ) ? ( n439 ) : ( x10 ) ;
assign n441 =  ( n424 ) ? ( n333 ) : ( x10 ) ;
assign n442 =  ( n424 ) ? ( n336 ) : ( x10 ) ;
assign n443 =  ( n424 ) ? ( n339 ) : ( x10 ) ;
assign n444 =  ( n424 ) ? ( n341 ) : ( x10 ) ;
assign n445 =  ( n424 ) ? ( n162 ) : ( x10 ) ;
assign n446 =  ( n424 ) ? ( n347 ) : ( x10 ) ;
assign n447 =  ( n424 ) ? ( n346 ) : ( x10 ) ;
assign n448 =  ( n424 ) ? ( n370 ) : ( x10 ) ;
assign n449 =  ( n424 ) ? ( n378 ) : ( x10 ) ;
assign n450 =  ( n424 ) ? ( n387 ) : ( x10 ) ;
assign n451 =  ( n424 ) ? ( n393 ) : ( x10 ) ;
assign n452 =  ( n424 ) ? ( n395 ) : ( x10 ) ;
assign n453 =  ( n230 ) ? ( n452 ) : ( x10 ) ;
assign n454 =  ( n229 ) ? ( n451 ) : ( n453 ) ;
assign n455 =  ( n228 ) ? ( n450 ) : ( n454 ) ;
assign n456 =  ( n227 ) ? ( n449 ) : ( n455 ) ;
assign n457 =  ( n226 ) ? ( n448 ) : ( n456 ) ;
assign n458 =  ( n220 ) ? ( n447 ) : ( n457 ) ;
assign n459 =  ( n219 ) ? ( n446 ) : ( n458 ) ;
assign n460 =  ( n343 ) ? ( n445 ) : ( n459 ) ;
assign n461 =  ( n218 ) ? ( n444 ) : ( n460 ) ;
assign n462 =  ( n217 ) ? ( n443 ) : ( n461 ) ;
assign n463 =  ( n216 ) ? ( n442 ) : ( n462 ) ;
assign n464 =  ( n215 ) ? ( n441 ) : ( n463 ) ;
assign n465 =  ( n214 ) ? ( n440 ) : ( n464 ) ;
assign n466 =  ( n213 ) ? ( n438 ) : ( n465 ) ;
assign n467 =  ( n212 ) ? ( n437 ) : ( n466 ) ;
assign n468 =  ( n210 ) ? ( n436 ) : ( n467 ) ;
assign n469 =  ( n209 ) ? ( n435 ) : ( n468 ) ;
assign n470 =  ( n206 ) ? ( n434 ) : ( n469 ) ;
assign n471 =  ( n205 ) ? ( n433 ) : ( n470 ) ;
assign n472 =  ( n202 ) ? ( n432 ) : ( n471 ) ;
assign n473 =  ( n199 ) ? ( n431 ) : ( n472 ) ;
assign n474 =  ( n197 ) ? ( n430 ) : ( n473 ) ;
assign n475 =  ( n195 ) ? ( n429 ) : ( n474 ) ;
assign n476 =  ( n193 ) ? ( n428 ) : ( n475 ) ;
assign n477 =  ( n191 ) ? ( n427 ) : ( n476 ) ;
assign n478 =  ( n189 ) ? ( n426 ) : ( n477 ) ;
assign n479 =  ( n187 ) ? ( n425 ) : ( n478 ) ;
assign n480 =  ( n296 ) == ( 5'd11 )  ;
assign n481 =  ( n480 ) ? ( n300 ) : ( x11 ) ;
assign n482 =  ( n480 ) ? ( n302 ) : ( x11 ) ;
assign n483 =  ( n480 ) ? ( n304 ) : ( x11 ) ;
assign n484 =  ( n480 ) ? ( n306 ) : ( x11 ) ;
assign n485 =  ( n480 ) ? ( n308 ) : ( x11 ) ;
assign n486 =  ( n480 ) ? ( n310 ) : ( x11 ) ;
assign n487 =  ( n480 ) ? ( n312 ) : ( x11 ) ;
assign n488 =  ( n480 ) ? ( n314 ) : ( x11 ) ;
assign n489 =  ( n480 ) ? ( n316 ) : ( x11 ) ;
assign n490 =  ( n480 ) ? ( n318 ) : ( x11 ) ;
assign n491 =  ( n480 ) ? ( n321 ) : ( x11 ) ;
assign n492 =  ( n480 ) ? ( n323 ) : ( x11 ) ;
assign n493 =  ( n480 ) ? ( n325 ) : ( x11 ) ;
assign n494 =  ( n480 ) ? ( n328 ) : ( x11 ) ;
assign n495 =  ( n480 ) ? ( n439 ) : ( x11 ) ;
assign n496 =  ( n480 ) ? ( n333 ) : ( x11 ) ;
assign n497 =  ( n480 ) ? ( n336 ) : ( x11 ) ;
assign n498 =  ( n480 ) ? ( n339 ) : ( x11 ) ;
assign n499 =  ( n480 ) ? ( n341 ) : ( x11 ) ;
assign n500 =  ( n480 ) ? ( n162 ) : ( x11 ) ;
assign n501 =  ( n480 ) ? ( n347 ) : ( x11 ) ;
assign n502 =  ( n480 ) ? ( n346 ) : ( x11 ) ;
assign n503 =  ( n480 ) ? ( n370 ) : ( x11 ) ;
assign n504 =  ( n480 ) ? ( n378 ) : ( x11 ) ;
assign n505 =  ( n480 ) ? ( n387 ) : ( x11 ) ;
assign n506 =  ( n480 ) ? ( n393 ) : ( x11 ) ;
assign n507 =  ( n480 ) ? ( n395 ) : ( x11 ) ;
assign n508 =  ( n230 ) ? ( n507 ) : ( x11 ) ;
assign n509 =  ( n229 ) ? ( n506 ) : ( n508 ) ;
assign n510 =  ( n228 ) ? ( n505 ) : ( n509 ) ;
assign n511 =  ( n227 ) ? ( n504 ) : ( n510 ) ;
assign n512 =  ( n226 ) ? ( n503 ) : ( n511 ) ;
assign n513 =  ( n220 ) ? ( n502 ) : ( n512 ) ;
assign n514 =  ( n219 ) ? ( n501 ) : ( n513 ) ;
assign n515 =  ( n343 ) ? ( n500 ) : ( n514 ) ;
assign n516 =  ( n218 ) ? ( n499 ) : ( n515 ) ;
assign n517 =  ( n217 ) ? ( n498 ) : ( n516 ) ;
assign n518 =  ( n216 ) ? ( n497 ) : ( n517 ) ;
assign n519 =  ( n215 ) ? ( n496 ) : ( n518 ) ;
assign n520 =  ( n214 ) ? ( n495 ) : ( n519 ) ;
assign n521 =  ( n213 ) ? ( n494 ) : ( n520 ) ;
assign n522 =  ( n212 ) ? ( n493 ) : ( n521 ) ;
assign n523 =  ( n210 ) ? ( n492 ) : ( n522 ) ;
assign n524 =  ( n209 ) ? ( n491 ) : ( n523 ) ;
assign n525 =  ( n206 ) ? ( n490 ) : ( n524 ) ;
assign n526 =  ( n205 ) ? ( n489 ) : ( n525 ) ;
assign n527 =  ( n202 ) ? ( n488 ) : ( n526 ) ;
assign n528 =  ( n199 ) ? ( n487 ) : ( n527 ) ;
assign n529 =  ( n197 ) ? ( n486 ) : ( n528 ) ;
assign n530 =  ( n195 ) ? ( n485 ) : ( n529 ) ;
assign n531 =  ( n193 ) ? ( n484 ) : ( n530 ) ;
assign n532 =  ( n191 ) ? ( n483 ) : ( n531 ) ;
assign n533 =  ( n189 ) ? ( n482 ) : ( n532 ) ;
assign n534 =  ( n187 ) ? ( n481 ) : ( n533 ) ;
assign n535 =  ( n296 ) == ( 5'd12 )  ;
assign n536 =  ( n535 ) ? ( n300 ) : ( x12 ) ;
assign n537 =  ( n535 ) ? ( n302 ) : ( x12 ) ;
assign n538 =  ( n535 ) ? ( n304 ) : ( x12 ) ;
assign n539 =  ( n535 ) ? ( n306 ) : ( x12 ) ;
assign n540 =  ( n535 ) ? ( n308 ) : ( x12 ) ;
assign n541 =  ( n535 ) ? ( n310 ) : ( x12 ) ;
assign n542 =  ( n535 ) ? ( n312 ) : ( x12 ) ;
assign n543 =  ( n535 ) ? ( n314 ) : ( x12 ) ;
assign n544 =  ( n535 ) ? ( n316 ) : ( x12 ) ;
assign n545 =  ( n535 ) ? ( n318 ) : ( x12 ) ;
assign n546 =  ( n535 ) ? ( n321 ) : ( x12 ) ;
assign n547 =  ( n535 ) ? ( n323 ) : ( x12 ) ;
assign n548 =  ( n535 ) ? ( n325 ) : ( x12 ) ;
assign n549 =  ( n535 ) ? ( n328 ) : ( x12 ) ;
assign n550 =  ( n535 ) ? ( n439 ) : ( x12 ) ;
assign n551 =  ( n535 ) ? ( n333 ) : ( x12 ) ;
assign n552 =  ( n70 ) < ( n327 )  ;
assign n553 =  ( n552 ) ? ( 32'd1 ) : ( 32'd0 ) ;
assign n554 =  ( n535 ) ? ( n553 ) : ( x12 ) ;
assign n555 =  ( n535 ) ? ( n339 ) : ( x12 ) ;
assign n556 =  ( n535 ) ? ( n341 ) : ( x12 ) ;
assign n557 =  ( n535 ) ? ( n162 ) : ( x12 ) ;
assign n558 =  ( n535 ) ? ( n347 ) : ( x12 ) ;
assign n559 =  ( n535 ) ? ( n346 ) : ( x12 ) ;
assign n560 =  ( n535 ) ? ( n370 ) : ( x12 ) ;
assign n561 =  ( n535 ) ? ( n378 ) : ( x12 ) ;
assign n562 =  ( n535 ) ? ( n387 ) : ( x12 ) ;
assign n563 =  ( n535 ) ? ( n393 ) : ( x12 ) ;
assign n564 =  ( n535 ) ? ( n395 ) : ( x12 ) ;
assign n565 =  ( n230 ) ? ( n564 ) : ( x12 ) ;
assign n566 =  ( n229 ) ? ( n563 ) : ( n565 ) ;
assign n567 =  ( n228 ) ? ( n562 ) : ( n566 ) ;
assign n568 =  ( n227 ) ? ( n561 ) : ( n567 ) ;
assign n569 =  ( n226 ) ? ( n560 ) : ( n568 ) ;
assign n570 =  ( n220 ) ? ( n559 ) : ( n569 ) ;
assign n571 =  ( n219 ) ? ( n558 ) : ( n570 ) ;
assign n572 =  ( n343 ) ? ( n557 ) : ( n571 ) ;
assign n573 =  ( n218 ) ? ( n556 ) : ( n572 ) ;
assign n574 =  ( n217 ) ? ( n555 ) : ( n573 ) ;
assign n575 =  ( n216 ) ? ( n554 ) : ( n574 ) ;
assign n576 =  ( n215 ) ? ( n551 ) : ( n575 ) ;
assign n577 =  ( n214 ) ? ( n550 ) : ( n576 ) ;
assign n578 =  ( n213 ) ? ( n549 ) : ( n577 ) ;
assign n579 =  ( n212 ) ? ( n548 ) : ( n578 ) ;
assign n580 =  ( n210 ) ? ( n547 ) : ( n579 ) ;
assign n581 =  ( n209 ) ? ( n546 ) : ( n580 ) ;
assign n582 =  ( n206 ) ? ( n545 ) : ( n581 ) ;
assign n583 =  ( n205 ) ? ( n544 ) : ( n582 ) ;
assign n584 =  ( n202 ) ? ( n543 ) : ( n583 ) ;
assign n585 =  ( n199 ) ? ( n542 ) : ( n584 ) ;
assign n586 =  ( n197 ) ? ( n541 ) : ( n585 ) ;
assign n587 =  ( n195 ) ? ( n540 ) : ( n586 ) ;
assign n588 =  ( n193 ) ? ( n539 ) : ( n587 ) ;
assign n589 =  ( n191 ) ? ( n538 ) : ( n588 ) ;
assign n590 =  ( n189 ) ? ( n537 ) : ( n589 ) ;
assign n591 =  ( n187 ) ? ( n536 ) : ( n590 ) ;
assign n592 =  ( n296 ) == ( 5'd13 )  ;
assign n593 =  ( n592 ) ? ( n300 ) : ( x13 ) ;
assign n594 =  ( n592 ) ? ( n302 ) : ( x13 ) ;
assign n595 =  ( n592 ) ? ( n304 ) : ( x13 ) ;
assign n596 =  ( n592 ) ? ( n306 ) : ( x13 ) ;
assign n597 =  ( n592 ) ? ( n308 ) : ( x13 ) ;
assign n598 =  ( n592 ) ? ( n310 ) : ( x13 ) ;
assign n599 =  ( n592 ) ? ( n312 ) : ( x13 ) ;
assign n600 =  ( n592 ) ? ( n314 ) : ( x13 ) ;
assign n601 =  ( n592 ) ? ( n316 ) : ( x13 ) ;
assign n602 =  ( n592 ) ? ( n318 ) : ( x13 ) ;
assign n603 =  ( n592 ) ? ( n321 ) : ( x13 ) ;
assign n604 =  ( n592 ) ? ( n323 ) : ( x13 ) ;
assign n605 =  ( n592 ) ? ( n325 ) : ( x13 ) ;
assign n606 =  ( n592 ) ? ( n328 ) : ( x13 ) ;
assign n607 =  ( n592 ) ? ( n439 ) : ( x13 ) ;
assign n608 =  ( n70 ) & ( n330 )  ;
assign n609 =  ( n592 ) ? ( n608 ) : ( x13 ) ;
assign n610 =  ( n592 ) ? ( n553 ) : ( x13 ) ;
assign n611 =  $signed( n70 ) < $signed( n330 )  ;
assign n612 =  ( n611 ) ? ( 32'd1 ) : ( 32'd0 ) ;
assign n613 =  ( n592 ) ? ( n612 ) : ( x13 ) ;
assign n614 =  ( n592 ) ? ( n341 ) : ( x13 ) ;
assign n615 =  ( n592 ) ? ( n162 ) : ( x13 ) ;
assign n616 =  ( n592 ) ? ( n347 ) : ( x13 ) ;
assign n617 =  ( n592 ) ? ( n346 ) : ( x13 ) ;
assign n618 =  ( n592 ) ? ( n370 ) : ( x13 ) ;
assign n619 =  ( n592 ) ? ( n378 ) : ( x13 ) ;
assign n620 =  ( n592 ) ? ( n387 ) : ( x13 ) ;
assign n621 =  ( n592 ) ? ( n393 ) : ( x13 ) ;
assign n622 =  ( n592 ) ? ( n395 ) : ( x13 ) ;
assign n623 =  ( n230 ) ? ( n622 ) : ( x13 ) ;
assign n624 =  ( n229 ) ? ( n621 ) : ( n623 ) ;
assign n625 =  ( n228 ) ? ( n620 ) : ( n624 ) ;
assign n626 =  ( n227 ) ? ( n619 ) : ( n625 ) ;
assign n627 =  ( n226 ) ? ( n618 ) : ( n626 ) ;
assign n628 =  ( n220 ) ? ( n617 ) : ( n627 ) ;
assign n629 =  ( n219 ) ? ( n616 ) : ( n628 ) ;
assign n630 =  ( n343 ) ? ( n615 ) : ( n629 ) ;
assign n631 =  ( n218 ) ? ( n614 ) : ( n630 ) ;
assign n632 =  ( n217 ) ? ( n613 ) : ( n631 ) ;
assign n633 =  ( n216 ) ? ( n610 ) : ( n632 ) ;
assign n634 =  ( n215 ) ? ( n609 ) : ( n633 ) ;
assign n635 =  ( n214 ) ? ( n607 ) : ( n634 ) ;
assign n636 =  ( n213 ) ? ( n606 ) : ( n635 ) ;
assign n637 =  ( n212 ) ? ( n605 ) : ( n636 ) ;
assign n638 =  ( n210 ) ? ( n604 ) : ( n637 ) ;
assign n639 =  ( n209 ) ? ( n603 ) : ( n638 ) ;
assign n640 =  ( n206 ) ? ( n602 ) : ( n639 ) ;
assign n641 =  ( n205 ) ? ( n601 ) : ( n640 ) ;
assign n642 =  ( n202 ) ? ( n600 ) : ( n641 ) ;
assign n643 =  ( n199 ) ? ( n599 ) : ( n642 ) ;
assign n644 =  ( n197 ) ? ( n598 ) : ( n643 ) ;
assign n645 =  ( n195 ) ? ( n597 ) : ( n644 ) ;
assign n646 =  ( n193 ) ? ( n596 ) : ( n645 ) ;
assign n647 =  ( n191 ) ? ( n595 ) : ( n646 ) ;
assign n648 =  ( n189 ) ? ( n594 ) : ( n647 ) ;
assign n649 =  ( n187 ) ? ( n593 ) : ( n648 ) ;
assign n650 =  ( n296 ) == ( 5'd14 )  ;
assign n651 =  ( n650 ) ? ( n300 ) : ( x14 ) ;
assign n652 =  ( n650 ) ? ( n302 ) : ( x14 ) ;
assign n653 =  ( n650 ) ? ( n304 ) : ( x14 ) ;
assign n654 =  ( n650 ) ? ( n306 ) : ( x14 ) ;
assign n655 =  ( n650 ) ? ( n308 ) : ( x14 ) ;
assign n656 =  ( n650 ) ? ( n310 ) : ( x14 ) ;
assign n657 =  ( n650 ) ? ( n312 ) : ( x14 ) ;
assign n658 =  ( n650 ) ? ( n314 ) : ( x14 ) ;
assign n659 =  ( n650 ) ? ( n316 ) : ( x14 ) ;
assign n660 =  ( n650 ) ? ( n318 ) : ( x14 ) ;
assign n661 =  ( n650 ) ? ( n321 ) : ( x14 ) ;
assign n662 =  ( n650 ) ? ( n323 ) : ( x14 ) ;
assign n663 =  ( n650 ) ? ( n325 ) : ( x14 ) ;
assign n664 =  ( n650 ) ? ( n328 ) : ( x14 ) ;
assign n665 =  ( n650 ) ? ( n439 ) : ( x14 ) ;
assign n666 =  ( n650 ) ? ( n333 ) : ( x14 ) ;
assign n667 =  ( n650 ) ? ( n553 ) : ( x14 ) ;
assign n668 =  ( n650 ) ? ( n339 ) : ( x14 ) ;
assign n669 =  ( n650 ) ? ( n341 ) : ( x14 ) ;
assign n670 =  ( n650 ) ? ( n162 ) : ( x14 ) ;
assign n671 =  ( n650 ) ? ( n347 ) : ( x14 ) ;
assign n672 =  ( n650 ) ? ( n346 ) : ( x14 ) ;
assign n673 =  ( n650 ) ? ( n370 ) : ( x14 ) ;
assign n674 =  ( n650 ) ? ( n378 ) : ( x14 ) ;
assign n675 =  ( n650 ) ? ( n387 ) : ( x14 ) ;
assign n676 =  ( n650 ) ? ( n393 ) : ( x14 ) ;
assign n677 =  ( n650 ) ? ( n395 ) : ( x14 ) ;
assign n678 =  ( n230 ) ? ( n677 ) : ( x14 ) ;
assign n679 =  ( n229 ) ? ( n676 ) : ( n678 ) ;
assign n680 =  ( n228 ) ? ( n675 ) : ( n679 ) ;
assign n681 =  ( n227 ) ? ( n674 ) : ( n680 ) ;
assign n682 =  ( n226 ) ? ( n673 ) : ( n681 ) ;
assign n683 =  ( n220 ) ? ( n672 ) : ( n682 ) ;
assign n684 =  ( n219 ) ? ( n671 ) : ( n683 ) ;
assign n685 =  ( n343 ) ? ( n670 ) : ( n684 ) ;
assign n686 =  ( n218 ) ? ( n669 ) : ( n685 ) ;
assign n687 =  ( n217 ) ? ( n668 ) : ( n686 ) ;
assign n688 =  ( n216 ) ? ( n667 ) : ( n687 ) ;
assign n689 =  ( n215 ) ? ( n666 ) : ( n688 ) ;
assign n690 =  ( n214 ) ? ( n665 ) : ( n689 ) ;
assign n691 =  ( n213 ) ? ( n664 ) : ( n690 ) ;
assign n692 =  ( n212 ) ? ( n663 ) : ( n691 ) ;
assign n693 =  ( n210 ) ? ( n662 ) : ( n692 ) ;
assign n694 =  ( n209 ) ? ( n661 ) : ( n693 ) ;
assign n695 =  ( n206 ) ? ( n660 ) : ( n694 ) ;
assign n696 =  ( n205 ) ? ( n659 ) : ( n695 ) ;
assign n697 =  ( n202 ) ? ( n658 ) : ( n696 ) ;
assign n698 =  ( n199 ) ? ( n657 ) : ( n697 ) ;
assign n699 =  ( n197 ) ? ( n656 ) : ( n698 ) ;
assign n700 =  ( n195 ) ? ( n655 ) : ( n699 ) ;
assign n701 =  ( n193 ) ? ( n654 ) : ( n700 ) ;
assign n702 =  ( n191 ) ? ( n653 ) : ( n701 ) ;
assign n703 =  ( n189 ) ? ( n652 ) : ( n702 ) ;
assign n704 =  ( n187 ) ? ( n651 ) : ( n703 ) ;
assign n705 =  ( n296 ) == ( 5'd15 )  ;
assign n706 =  ( n705 ) ? ( n300 ) : ( x15 ) ;
assign n707 =  ( n705 ) ? ( n302 ) : ( x15 ) ;
assign n708 =  ( n705 ) ? ( n304 ) : ( x15 ) ;
assign n709 =  ( n705 ) ? ( n306 ) : ( x15 ) ;
assign n710 =  ( n705 ) ? ( n308 ) : ( x15 ) ;
assign n711 =  ( n705 ) ? ( n310 ) : ( x15 ) ;
assign n712 =  ( n705 ) ? ( n312 ) : ( x15 ) ;
assign n713 =  ( n705 ) ? ( n314 ) : ( x15 ) ;
assign n714 =  ( n705 ) ? ( n316 ) : ( x15 ) ;
assign n715 =  ( n705 ) ? ( n318 ) : ( x15 ) ;
assign n716 =  ( n705 ) ? ( n321 ) : ( x15 ) ;
assign n717 =  ( n705 ) ? ( n323 ) : ( x15 ) ;
assign n718 =  ( n705 ) ? ( n325 ) : ( x15 ) ;
assign n719 =  ( n70 ) ^ ( n330 )  ;
assign n720 =  ( n705 ) ? ( n719 ) : ( x15 ) ;
assign n721 =  ( n705 ) ? ( n439 ) : ( x15 ) ;
assign n722 =  ( n705 ) ? ( n333 ) : ( x15 ) ;
assign n723 =  ( n705 ) ? ( n336 ) : ( x15 ) ;
assign n724 =  ( n705 ) ? ( n339 ) : ( x15 ) ;
assign n725 =  ( n705 ) ? ( n341 ) : ( x15 ) ;
assign n726 =  ( n705 ) ? ( n162 ) : ( x15 ) ;
assign n727 =  ( n705 ) ? ( n347 ) : ( x15 ) ;
assign n728 =  ( n705 ) ? ( n346 ) : ( x15 ) ;
assign n729 =  ( n705 ) ? ( n370 ) : ( x15 ) ;
assign n730 =  ( n705 ) ? ( n378 ) : ( x15 ) ;
assign n731 =  ( n705 ) ? ( n387 ) : ( x15 ) ;
assign n732 =  ( n705 ) ? ( n393 ) : ( x15 ) ;
assign n733 =  ( n705 ) ? ( n395 ) : ( x15 ) ;
assign n734 =  ( n230 ) ? ( n733 ) : ( x15 ) ;
assign n735 =  ( n229 ) ? ( n732 ) : ( n734 ) ;
assign n736 =  ( n228 ) ? ( n731 ) : ( n735 ) ;
assign n737 =  ( n227 ) ? ( n730 ) : ( n736 ) ;
assign n738 =  ( n226 ) ? ( n729 ) : ( n737 ) ;
assign n739 =  ( n220 ) ? ( n728 ) : ( n738 ) ;
assign n740 =  ( n219 ) ? ( n727 ) : ( n739 ) ;
assign n741 =  ( n343 ) ? ( n726 ) : ( n740 ) ;
assign n742 =  ( n218 ) ? ( n725 ) : ( n741 ) ;
assign n743 =  ( n217 ) ? ( n724 ) : ( n742 ) ;
assign n744 =  ( n216 ) ? ( n723 ) : ( n743 ) ;
assign n745 =  ( n215 ) ? ( n722 ) : ( n744 ) ;
assign n746 =  ( n214 ) ? ( n721 ) : ( n745 ) ;
assign n747 =  ( n213 ) ? ( n720 ) : ( n746 ) ;
assign n748 =  ( n212 ) ? ( n718 ) : ( n747 ) ;
assign n749 =  ( n210 ) ? ( n717 ) : ( n748 ) ;
assign n750 =  ( n209 ) ? ( n716 ) : ( n749 ) ;
assign n751 =  ( n206 ) ? ( n715 ) : ( n750 ) ;
assign n752 =  ( n205 ) ? ( n714 ) : ( n751 ) ;
assign n753 =  ( n202 ) ? ( n713 ) : ( n752 ) ;
assign n754 =  ( n199 ) ? ( n712 ) : ( n753 ) ;
assign n755 =  ( n197 ) ? ( n711 ) : ( n754 ) ;
assign n756 =  ( n195 ) ? ( n710 ) : ( n755 ) ;
assign n757 =  ( n193 ) ? ( n709 ) : ( n756 ) ;
assign n758 =  ( n191 ) ? ( n708 ) : ( n757 ) ;
assign n759 =  ( n189 ) ? ( n707 ) : ( n758 ) ;
assign n760 =  ( n187 ) ? ( n706 ) : ( n759 ) ;
assign n761 =  ( n296 ) == ( 5'd16 )  ;
assign n762 =  ( n761 ) ? ( n300 ) : ( x16 ) ;
assign n763 =  ( n761 ) ? ( n302 ) : ( x16 ) ;
assign n764 =  ( n761 ) ? ( n304 ) : ( x16 ) ;
assign n765 =  ( n761 ) ? ( n306 ) : ( x16 ) ;
assign n766 =  ( n761 ) ? ( n308 ) : ( x16 ) ;
assign n767 =  ( n761 ) ? ( n310 ) : ( x16 ) ;
assign n768 =  ( n761 ) ? ( n312 ) : ( x16 ) ;
assign n769 =  ( n761 ) ? ( n314 ) : ( x16 ) ;
assign n770 =  ( n761 ) ? ( n316 ) : ( x16 ) ;
assign n771 =  ( n761 ) ? ( n318 ) : ( x16 ) ;
assign n772 =  ( n761 ) ? ( n321 ) : ( x16 ) ;
assign n773 =  ( n761 ) ? ( n323 ) : ( x16 ) ;
assign n774 =  ( n761 ) ? ( n325 ) : ( x16 ) ;
assign n775 =  ( n761 ) ? ( n328 ) : ( x16 ) ;
assign n776 =  ( n761 ) ? ( n439 ) : ( x16 ) ;
assign n777 =  ( n761 ) ? ( n333 ) : ( x16 ) ;
assign n778 =  ( n761 ) ? ( n553 ) : ( x16 ) ;
assign n779 =  ( n761 ) ? ( n339 ) : ( x16 ) ;
assign n780 =  ( n761 ) ? ( n341 ) : ( x16 ) ;
assign n781 =  ( n761 ) ? ( n162 ) : ( x16 ) ;
assign n782 =  ( n761 ) ? ( n347 ) : ( x16 ) ;
assign n783 =  ( n761 ) ? ( n346 ) : ( x16 ) ;
assign n784 =  ( n761 ) ? ( n370 ) : ( x16 ) ;
assign n785 =  ( n761 ) ? ( n378 ) : ( x16 ) ;
assign n786 =  ( n761 ) ? ( n387 ) : ( x16 ) ;
assign n787 =  ( n761 ) ? ( n393 ) : ( x16 ) ;
assign n788 =  ( n761 ) ? ( n395 ) : ( x16 ) ;
assign n789 =  ( n230 ) ? ( n788 ) : ( x16 ) ;
assign n790 =  ( n229 ) ? ( n787 ) : ( n789 ) ;
assign n791 =  ( n228 ) ? ( n786 ) : ( n790 ) ;
assign n792 =  ( n227 ) ? ( n785 ) : ( n791 ) ;
assign n793 =  ( n226 ) ? ( n784 ) : ( n792 ) ;
assign n794 =  ( n220 ) ? ( n783 ) : ( n793 ) ;
assign n795 =  ( n219 ) ? ( n782 ) : ( n794 ) ;
assign n796 =  ( n343 ) ? ( n781 ) : ( n795 ) ;
assign n797 =  ( n218 ) ? ( n780 ) : ( n796 ) ;
assign n798 =  ( n217 ) ? ( n779 ) : ( n797 ) ;
assign n799 =  ( n216 ) ? ( n778 ) : ( n798 ) ;
assign n800 =  ( n215 ) ? ( n777 ) : ( n799 ) ;
assign n801 =  ( n214 ) ? ( n776 ) : ( n800 ) ;
assign n802 =  ( n213 ) ? ( n775 ) : ( n801 ) ;
assign n803 =  ( n212 ) ? ( n774 ) : ( n802 ) ;
assign n804 =  ( n210 ) ? ( n773 ) : ( n803 ) ;
assign n805 =  ( n209 ) ? ( n772 ) : ( n804 ) ;
assign n806 =  ( n206 ) ? ( n771 ) : ( n805 ) ;
assign n807 =  ( n205 ) ? ( n770 ) : ( n806 ) ;
assign n808 =  ( n202 ) ? ( n769 ) : ( n807 ) ;
assign n809 =  ( n199 ) ? ( n768 ) : ( n808 ) ;
assign n810 =  ( n197 ) ? ( n767 ) : ( n809 ) ;
assign n811 =  ( n195 ) ? ( n766 ) : ( n810 ) ;
assign n812 =  ( n193 ) ? ( n765 ) : ( n811 ) ;
assign n813 =  ( n191 ) ? ( n764 ) : ( n812 ) ;
assign n814 =  ( n189 ) ? ( n763 ) : ( n813 ) ;
assign n815 =  ( n187 ) ? ( n762 ) : ( n814 ) ;
assign n816 =  ( n296 ) == ( 5'd17 )  ;
assign n817 =  ( n816 ) ? ( n300 ) : ( x17 ) ;
assign n818 =  ( n816 ) ? ( n302 ) : ( x17 ) ;
assign n819 =  ( n816 ) ? ( n304 ) : ( x17 ) ;
assign n820 =  ( n816 ) ? ( n306 ) : ( x17 ) ;
assign n821 =  ( n816 ) ? ( n308 ) : ( x17 ) ;
assign n822 =  ( n816 ) ? ( n310 ) : ( x17 ) ;
assign n823 =  ( n816 ) ? ( n312 ) : ( x17 ) ;
assign n824 =  ( n816 ) ? ( n314 ) : ( x17 ) ;
assign n825 =  ( n816 ) ? ( n316 ) : ( x17 ) ;
assign n826 =  ( n816 ) ? ( n318 ) : ( x17 ) ;
assign n827 =  ( n816 ) ? ( n321 ) : ( x17 ) ;
assign n828 =  ( n816 ) ? ( n323 ) : ( x17 ) ;
assign n829 =  ( n816 ) ? ( n325 ) : ( x17 ) ;
assign n830 =  ( n816 ) ? ( n328 ) : ( x17 ) ;
assign n831 =  ( n816 ) ? ( n439 ) : ( x17 ) ;
assign n832 =  ( n816 ) ? ( n333 ) : ( x17 ) ;
assign n833 =  ( n816 ) ? ( n553 ) : ( x17 ) ;
assign n834 =  ( n816 ) ? ( n339 ) : ( x17 ) ;
assign n835 =  ( n816 ) ? ( n341 ) : ( x17 ) ;
assign n836 =  ( n816 ) ? ( n162 ) : ( x17 ) ;
assign n837 =  ( n816 ) ? ( n347 ) : ( x17 ) ;
assign n838 =  ( n816 ) ? ( n346 ) : ( x17 ) ;
assign n839 =  ( n816 ) ? ( n370 ) : ( x17 ) ;
assign n840 =  ( n816 ) ? ( n378 ) : ( x17 ) ;
assign n841 =  ( n816 ) ? ( n387 ) : ( x17 ) ;
assign n842 =  ( n816 ) ? ( n393 ) : ( x17 ) ;
assign n843 =  ( n816 ) ? ( n395 ) : ( x17 ) ;
assign n844 =  ( n230 ) ? ( n843 ) : ( x17 ) ;
assign n845 =  ( n229 ) ? ( n842 ) : ( n844 ) ;
assign n846 =  ( n228 ) ? ( n841 ) : ( n845 ) ;
assign n847 =  ( n227 ) ? ( n840 ) : ( n846 ) ;
assign n848 =  ( n226 ) ? ( n839 ) : ( n847 ) ;
assign n849 =  ( n220 ) ? ( n838 ) : ( n848 ) ;
assign n850 =  ( n219 ) ? ( n837 ) : ( n849 ) ;
assign n851 =  ( n343 ) ? ( n836 ) : ( n850 ) ;
assign n852 =  ( n218 ) ? ( n835 ) : ( n851 ) ;
assign n853 =  ( n217 ) ? ( n834 ) : ( n852 ) ;
assign n854 =  ( n216 ) ? ( n833 ) : ( n853 ) ;
assign n855 =  ( n215 ) ? ( n832 ) : ( n854 ) ;
assign n856 =  ( n214 ) ? ( n831 ) : ( n855 ) ;
assign n857 =  ( n213 ) ? ( n830 ) : ( n856 ) ;
assign n858 =  ( n212 ) ? ( n829 ) : ( n857 ) ;
assign n859 =  ( n210 ) ? ( n828 ) : ( n858 ) ;
assign n860 =  ( n209 ) ? ( n827 ) : ( n859 ) ;
assign n861 =  ( n206 ) ? ( n826 ) : ( n860 ) ;
assign n862 =  ( n205 ) ? ( n825 ) : ( n861 ) ;
assign n863 =  ( n202 ) ? ( n824 ) : ( n862 ) ;
assign n864 =  ( n199 ) ? ( n823 ) : ( n863 ) ;
assign n865 =  ( n197 ) ? ( n822 ) : ( n864 ) ;
assign n866 =  ( n195 ) ? ( n821 ) : ( n865 ) ;
assign n867 =  ( n193 ) ? ( n820 ) : ( n866 ) ;
assign n868 =  ( n191 ) ? ( n819 ) : ( n867 ) ;
assign n869 =  ( n189 ) ? ( n818 ) : ( n868 ) ;
assign n870 =  ( n187 ) ? ( n817 ) : ( n869 ) ;
assign n871 =  ( n296 ) == ( 5'd18 )  ;
assign n872 =  ( n871 ) ? ( n300 ) : ( x18 ) ;
assign n873 =  ( n871 ) ? ( n302 ) : ( x18 ) ;
assign n874 =  ( n871 ) ? ( n304 ) : ( x18 ) ;
assign n875 =  ( n871 ) ? ( n306 ) : ( x18 ) ;
assign n876 =  ( n871 ) ? ( n308 ) : ( x18 ) ;
assign n877 =  ( n871 ) ? ( n310 ) : ( x18 ) ;
assign n878 =  ( n871 ) ? ( n312 ) : ( x18 ) ;
assign n879 =  ( n871 ) ? ( n314 ) : ( x18 ) ;
assign n880 =  ( n871 ) ? ( n316 ) : ( x18 ) ;
assign n881 =  ( n871 ) ? ( n318 ) : ( x18 ) ;
assign n882 =  ( n871 ) ? ( n321 ) : ( x18 ) ;
assign n883 =  ( n871 ) ? ( n323 ) : ( x18 ) ;
assign n884 =  ( n871 ) ? ( n325 ) : ( x18 ) ;
assign n885 =  ( n871 ) ? ( n328 ) : ( x18 ) ;
assign n886 =  ( n871 ) ? ( n439 ) : ( x18 ) ;
assign n887 =  ( n871 ) ? ( n608 ) : ( x18 ) ;
assign n888 =  ( n871 ) ? ( n553 ) : ( x18 ) ;
assign n889 =  ( n871 ) ? ( n339 ) : ( x18 ) ;
assign n890 =  ( n871 ) ? ( n341 ) : ( x18 ) ;
assign n891 =  ( n871 ) ? ( n162 ) : ( x18 ) ;
assign n892 =  ( n871 ) ? ( n347 ) : ( x18 ) ;
assign n893 =  ( n871 ) ? ( n346 ) : ( x18 ) ;
assign n894 =  ( n871 ) ? ( n370 ) : ( x18 ) ;
assign n895 =  ( n871 ) ? ( n378 ) : ( x18 ) ;
assign n896 =  ( n871 ) ? ( n387 ) : ( x18 ) ;
assign n897 =  ( n871 ) ? ( n393 ) : ( x18 ) ;
assign n898 =  ( n871 ) ? ( n395 ) : ( x18 ) ;
assign n899 =  ( n230 ) ? ( n898 ) : ( x18 ) ;
assign n900 =  ( n229 ) ? ( n897 ) : ( n899 ) ;
assign n901 =  ( n228 ) ? ( n896 ) : ( n900 ) ;
assign n902 =  ( n227 ) ? ( n895 ) : ( n901 ) ;
assign n903 =  ( n226 ) ? ( n894 ) : ( n902 ) ;
assign n904 =  ( n220 ) ? ( n893 ) : ( n903 ) ;
assign n905 =  ( n219 ) ? ( n892 ) : ( n904 ) ;
assign n906 =  ( n343 ) ? ( n891 ) : ( n905 ) ;
assign n907 =  ( n218 ) ? ( n890 ) : ( n906 ) ;
assign n908 =  ( n217 ) ? ( n889 ) : ( n907 ) ;
assign n909 =  ( n216 ) ? ( n888 ) : ( n908 ) ;
assign n910 =  ( n215 ) ? ( n887 ) : ( n909 ) ;
assign n911 =  ( n214 ) ? ( n886 ) : ( n910 ) ;
assign n912 =  ( n213 ) ? ( n885 ) : ( n911 ) ;
assign n913 =  ( n212 ) ? ( n884 ) : ( n912 ) ;
assign n914 =  ( n210 ) ? ( n883 ) : ( n913 ) ;
assign n915 =  ( n209 ) ? ( n882 ) : ( n914 ) ;
assign n916 =  ( n206 ) ? ( n881 ) : ( n915 ) ;
assign n917 =  ( n205 ) ? ( n880 ) : ( n916 ) ;
assign n918 =  ( n202 ) ? ( n879 ) : ( n917 ) ;
assign n919 =  ( n199 ) ? ( n878 ) : ( n918 ) ;
assign n920 =  ( n197 ) ? ( n877 ) : ( n919 ) ;
assign n921 =  ( n195 ) ? ( n876 ) : ( n920 ) ;
assign n922 =  ( n193 ) ? ( n875 ) : ( n921 ) ;
assign n923 =  ( n191 ) ? ( n874 ) : ( n922 ) ;
assign n924 =  ( n189 ) ? ( n873 ) : ( n923 ) ;
assign n925 =  ( n187 ) ? ( n872 ) : ( n924 ) ;
assign n926 =  ( n296 ) == ( 5'd19 )  ;
assign n927 =  ( n926 ) ? ( n300 ) : ( x19 ) ;
assign n928 =  ( n926 ) ? ( n302 ) : ( x19 ) ;
assign n929 =  ( n926 ) ? ( n304 ) : ( x19 ) ;
assign n930 =  ( n926 ) ? ( n306 ) : ( x19 ) ;
assign n931 =  ( n926 ) ? ( n308 ) : ( x19 ) ;
assign n932 =  ( n926 ) ? ( n310 ) : ( x19 ) ;
assign n933 =  ( n926 ) ? ( n312 ) : ( x19 ) ;
assign n934 =  ( n926 ) ? ( n314 ) : ( x19 ) ;
assign n935 =  ( n926 ) ? ( n316 ) : ( x19 ) ;
assign n936 =  ( n926 ) ? ( n318 ) : ( x19 ) ;
assign n937 =  ( n926 ) ? ( n321 ) : ( x19 ) ;
assign n938 =  ( n926 ) ? ( n323 ) : ( x19 ) ;
assign n939 =  ( n926 ) ? ( n325 ) : ( x19 ) ;
assign n940 =  ( n926 ) ? ( n328 ) : ( x19 ) ;
assign n941 =  ( n926 ) ? ( n331 ) : ( x19 ) ;
assign n942 =  ( n926 ) ? ( n333 ) : ( x19 ) ;
assign n943 =  ( n926 ) ? ( n553 ) : ( x19 ) ;
assign n944 =  ( n926 ) ? ( n339 ) : ( x19 ) ;
assign n945 =  ( n926 ) ? ( n341 ) : ( x19 ) ;
assign n946 =  ( n926 ) ? ( n162 ) : ( x19 ) ;
assign n947 =  ( n926 ) ? ( n347 ) : ( x19 ) ;
assign n948 =  ( n926 ) ? ( n346 ) : ( x19 ) ;
assign n949 =  ( n926 ) ? ( n370 ) : ( x19 ) ;
assign n950 =  ( n926 ) ? ( n378 ) : ( x19 ) ;
assign n951 =  ( n926 ) ? ( n387 ) : ( x19 ) ;
assign n952 =  ( n926 ) ? ( n393 ) : ( x19 ) ;
assign n953 =  ( n926 ) ? ( n395 ) : ( x19 ) ;
assign n954 =  ( n230 ) ? ( n953 ) : ( x19 ) ;
assign n955 =  ( n229 ) ? ( n952 ) : ( n954 ) ;
assign n956 =  ( n228 ) ? ( n951 ) : ( n955 ) ;
assign n957 =  ( n227 ) ? ( n950 ) : ( n956 ) ;
assign n958 =  ( n226 ) ? ( n949 ) : ( n957 ) ;
assign n959 =  ( n220 ) ? ( n948 ) : ( n958 ) ;
assign n960 =  ( n219 ) ? ( n947 ) : ( n959 ) ;
assign n961 =  ( n343 ) ? ( n946 ) : ( n960 ) ;
assign n962 =  ( n218 ) ? ( n945 ) : ( n961 ) ;
assign n963 =  ( n217 ) ? ( n944 ) : ( n962 ) ;
assign n964 =  ( n216 ) ? ( n943 ) : ( n963 ) ;
assign n965 =  ( n215 ) ? ( n942 ) : ( n964 ) ;
assign n966 =  ( n214 ) ? ( n941 ) : ( n965 ) ;
assign n967 =  ( n213 ) ? ( n940 ) : ( n966 ) ;
assign n968 =  ( n212 ) ? ( n939 ) : ( n967 ) ;
assign n969 =  ( n210 ) ? ( n938 ) : ( n968 ) ;
assign n970 =  ( n209 ) ? ( n937 ) : ( n969 ) ;
assign n971 =  ( n206 ) ? ( n936 ) : ( n970 ) ;
assign n972 =  ( n205 ) ? ( n935 ) : ( n971 ) ;
assign n973 =  ( n202 ) ? ( n934 ) : ( n972 ) ;
assign n974 =  ( n199 ) ? ( n933 ) : ( n973 ) ;
assign n975 =  ( n197 ) ? ( n932 ) : ( n974 ) ;
assign n976 =  ( n195 ) ? ( n931 ) : ( n975 ) ;
assign n977 =  ( n193 ) ? ( n930 ) : ( n976 ) ;
assign n978 =  ( n191 ) ? ( n929 ) : ( n977 ) ;
assign n979 =  ( n189 ) ? ( n928 ) : ( n978 ) ;
assign n980 =  ( n187 ) ? ( n927 ) : ( n979 ) ;
assign n981 =  ( n296 ) == ( 5'd2 )  ;
assign n982 =  ( n981 ) ? ( n300 ) : ( x2 ) ;
assign n983 =  ( n981 ) ? ( n302 ) : ( x2 ) ;
assign n984 =  ( n981 ) ? ( n304 ) : ( x2 ) ;
assign n985 =  ( n981 ) ? ( n306 ) : ( x2 ) ;
assign n986 =  ( n981 ) ? ( n308 ) : ( x2 ) ;
assign n987 =  ( n981 ) ? ( n310 ) : ( x2 ) ;
assign n988 =  ( n981 ) ? ( n312 ) : ( x2 ) ;
assign n989 =  ( n981 ) ? ( n314 ) : ( x2 ) ;
assign n990 =  ( n981 ) ? ( n316 ) : ( x2 ) ;
assign n991 =  ( n981 ) ? ( n318 ) : ( x2 ) ;
assign n992 =  ( n981 ) ? ( n321 ) : ( x2 ) ;
assign n993 =  ( n981 ) ? ( n323 ) : ( x2 ) ;
assign n994 =  ( n981 ) ? ( n325 ) : ( x2 ) ;
assign n995 =  ( n981 ) ? ( n328 ) : ( x2 ) ;
assign n996 =  ( n981 ) ? ( n439 ) : ( x2 ) ;
assign n997 =  ( n981 ) ? ( n333 ) : ( x2 ) ;
assign n998 =  ( n981 ) ? ( n553 ) : ( x2 ) ;
assign n999 =  ( n981 ) ? ( n339 ) : ( x2 ) ;
assign n1000 =  ( n981 ) ? ( n341 ) : ( x2 ) ;
assign n1001 =  ( n981 ) ? ( n162 ) : ( x2 ) ;
assign n1002 =  ( n981 ) ? ( n347 ) : ( x2 ) ;
assign n1003 =  ( n981 ) ? ( n346 ) : ( x2 ) ;
assign n1004 =  ( n981 ) ? ( n370 ) : ( x2 ) ;
assign n1005 =  ( n981 ) ? ( n378 ) : ( x2 ) ;
assign n1006 =  ( n981 ) ? ( n387 ) : ( x2 ) ;
assign n1007 =  ( n981 ) ? ( n393 ) : ( x2 ) ;
assign n1008 =  ( n981 ) ? ( n395 ) : ( x2 ) ;
assign n1009 =  ( n230 ) ? ( n1008 ) : ( x2 ) ;
assign n1010 =  ( n229 ) ? ( n1007 ) : ( n1009 ) ;
assign n1011 =  ( n228 ) ? ( n1006 ) : ( n1010 ) ;
assign n1012 =  ( n227 ) ? ( n1005 ) : ( n1011 ) ;
assign n1013 =  ( n226 ) ? ( n1004 ) : ( n1012 ) ;
assign n1014 =  ( n220 ) ? ( n1003 ) : ( n1013 ) ;
assign n1015 =  ( n219 ) ? ( n1002 ) : ( n1014 ) ;
assign n1016 =  ( n343 ) ? ( n1001 ) : ( n1015 ) ;
assign n1017 =  ( n218 ) ? ( n1000 ) : ( n1016 ) ;
assign n1018 =  ( n217 ) ? ( n999 ) : ( n1017 ) ;
assign n1019 =  ( n216 ) ? ( n998 ) : ( n1018 ) ;
assign n1020 =  ( n215 ) ? ( n997 ) : ( n1019 ) ;
assign n1021 =  ( n214 ) ? ( n996 ) : ( n1020 ) ;
assign n1022 =  ( n213 ) ? ( n995 ) : ( n1021 ) ;
assign n1023 =  ( n212 ) ? ( n994 ) : ( n1022 ) ;
assign n1024 =  ( n210 ) ? ( n993 ) : ( n1023 ) ;
assign n1025 =  ( n209 ) ? ( n992 ) : ( n1024 ) ;
assign n1026 =  ( n206 ) ? ( n991 ) : ( n1025 ) ;
assign n1027 =  ( n205 ) ? ( n990 ) : ( n1026 ) ;
assign n1028 =  ( n202 ) ? ( n989 ) : ( n1027 ) ;
assign n1029 =  ( n199 ) ? ( n988 ) : ( n1028 ) ;
assign n1030 =  ( n197 ) ? ( n987 ) : ( n1029 ) ;
assign n1031 =  ( n195 ) ? ( n986 ) : ( n1030 ) ;
assign n1032 =  ( n193 ) ? ( n985 ) : ( n1031 ) ;
assign n1033 =  ( n191 ) ? ( n984 ) : ( n1032 ) ;
assign n1034 =  ( n189 ) ? ( n983 ) : ( n1033 ) ;
assign n1035 =  ( n187 ) ? ( n982 ) : ( n1034 ) ;
assign n1036 =  ( n296 ) == ( 5'd20 )  ;
assign n1037 =  ( n1036 ) ? ( n300 ) : ( x20 ) ;
assign n1038 =  ( n1036 ) ? ( n302 ) : ( x20 ) ;
assign n1039 =  ( n1036 ) ? ( n304 ) : ( x20 ) ;
assign n1040 =  ( n1036 ) ? ( n306 ) : ( x20 ) ;
assign n1041 =  ( n1036 ) ? ( n308 ) : ( x20 ) ;
assign n1042 =  ( n1036 ) ? ( n310 ) : ( x20 ) ;
assign n1043 =  ( n1036 ) ? ( n312 ) : ( x20 ) ;
assign n1044 =  ( n1036 ) ? ( n314 ) : ( x20 ) ;
assign n1045 =  ( n1036 ) ? ( n316 ) : ( x20 ) ;
assign n1046 =  ( n1036 ) ? ( n318 ) : ( x20 ) ;
assign n1047 =  ( n1036 ) ? ( n321 ) : ( x20 ) ;
assign n1048 =  ( n1036 ) ? ( n323 ) : ( x20 ) ;
assign n1049 =  ( n1036 ) ? ( n325 ) : ( x20 ) ;
assign n1050 =  ( n1036 ) ? ( n328 ) : ( x20 ) ;
assign n1051 =  ( n1036 ) ? ( n439 ) : ( x20 ) ;
assign n1052 =  ( n1036 ) ? ( n333 ) : ( x20 ) ;
assign n1053 =  ( n1036 ) ? ( n336 ) : ( x20 ) ;
assign n1054 =  ( n1036 ) ? ( n339 ) : ( x20 ) ;
assign n1055 =  ( n1036 ) ? ( n341 ) : ( x20 ) ;
assign n1056 =  ( n1036 ) ? ( n162 ) : ( x20 ) ;
assign n1057 =  ( n1036 ) ? ( n347 ) : ( x20 ) ;
assign n1058 =  ( n1036 ) ? ( n346 ) : ( x20 ) ;
assign n1059 =  ( n1036 ) ? ( n370 ) : ( x20 ) ;
assign n1060 =  ( n1036 ) ? ( n378 ) : ( x20 ) ;
assign n1061 =  ( n1036 ) ? ( n387 ) : ( x20 ) ;
assign n1062 =  ( n1036 ) ? ( n393 ) : ( x20 ) ;
assign n1063 =  ( n1036 ) ? ( n395 ) : ( x20 ) ;
assign n1064 =  ( n230 ) ? ( n1063 ) : ( x20 ) ;
assign n1065 =  ( n229 ) ? ( n1062 ) : ( n1064 ) ;
assign n1066 =  ( n228 ) ? ( n1061 ) : ( n1065 ) ;
assign n1067 =  ( n227 ) ? ( n1060 ) : ( n1066 ) ;
assign n1068 =  ( n226 ) ? ( n1059 ) : ( n1067 ) ;
assign n1069 =  ( n220 ) ? ( n1058 ) : ( n1068 ) ;
assign n1070 =  ( n219 ) ? ( n1057 ) : ( n1069 ) ;
assign n1071 =  ( n343 ) ? ( n1056 ) : ( n1070 ) ;
assign n1072 =  ( n218 ) ? ( n1055 ) : ( n1071 ) ;
assign n1073 =  ( n217 ) ? ( n1054 ) : ( n1072 ) ;
assign n1074 =  ( n216 ) ? ( n1053 ) : ( n1073 ) ;
assign n1075 =  ( n215 ) ? ( n1052 ) : ( n1074 ) ;
assign n1076 =  ( n214 ) ? ( n1051 ) : ( n1075 ) ;
assign n1077 =  ( n213 ) ? ( n1050 ) : ( n1076 ) ;
assign n1078 =  ( n212 ) ? ( n1049 ) : ( n1077 ) ;
assign n1079 =  ( n210 ) ? ( n1048 ) : ( n1078 ) ;
assign n1080 =  ( n209 ) ? ( n1047 ) : ( n1079 ) ;
assign n1081 =  ( n206 ) ? ( n1046 ) : ( n1080 ) ;
assign n1082 =  ( n205 ) ? ( n1045 ) : ( n1081 ) ;
assign n1083 =  ( n202 ) ? ( n1044 ) : ( n1082 ) ;
assign n1084 =  ( n199 ) ? ( n1043 ) : ( n1083 ) ;
assign n1085 =  ( n197 ) ? ( n1042 ) : ( n1084 ) ;
assign n1086 =  ( n195 ) ? ( n1041 ) : ( n1085 ) ;
assign n1087 =  ( n193 ) ? ( n1040 ) : ( n1086 ) ;
assign n1088 =  ( n191 ) ? ( n1039 ) : ( n1087 ) ;
assign n1089 =  ( n189 ) ? ( n1038 ) : ( n1088 ) ;
assign n1090 =  ( n187 ) ? ( n1037 ) : ( n1089 ) ;
assign n1091 =  ( n296 ) == ( 5'd21 )  ;
assign n1092 =  ( n1091 ) ? ( n300 ) : ( x21 ) ;
assign n1093 =  ( n1091 ) ? ( n302 ) : ( x21 ) ;
assign n1094 =  ( n1091 ) ? ( n304 ) : ( x21 ) ;
assign n1095 =  ( n1091 ) ? ( n306 ) : ( x21 ) ;
assign n1096 =  ( n1091 ) ? ( n308 ) : ( x21 ) ;
assign n1097 =  ( n1091 ) ? ( n310 ) : ( x21 ) ;
assign n1098 =  ( n1091 ) ? ( n312 ) : ( x21 ) ;
assign n1099 =  ( n1091 ) ? ( n314 ) : ( x21 ) ;
assign n1100 =  ( n1091 ) ? ( n316 ) : ( x21 ) ;
assign n1101 =  ( n1091 ) ? ( n318 ) : ( x21 ) ;
assign n1102 =  ( n1091 ) ? ( n321 ) : ( x21 ) ;
assign n1103 =  ( n1091 ) ? ( n323 ) : ( x21 ) ;
assign n1104 =  ( n1091 ) ? ( n325 ) : ( x21 ) ;
assign n1105 =  ( n1091 ) ? ( n328 ) : ( x21 ) ;
assign n1106 =  ( n1091 ) ? ( n439 ) : ( x21 ) ;
assign n1107 =  ( n1091 ) ? ( n608 ) : ( x21 ) ;
assign n1108 =  ( n1091 ) ? ( n553 ) : ( x21 ) ;
assign n1109 =  ( n1091 ) ? ( n612 ) : ( x21 ) ;
assign n1110 =  ( n1091 ) ? ( n341 ) : ( x21 ) ;
assign n1111 =  ( n1091 ) ? ( n162 ) : ( x21 ) ;
assign n1112 =  ( n1091 ) ? ( n347 ) : ( x21 ) ;
assign n1113 =  ( n1091 ) ? ( n346 ) : ( x21 ) ;
assign n1114 =  ( n1091 ) ? ( n370 ) : ( x21 ) ;
assign n1115 =  ( n1091 ) ? ( n378 ) : ( x21 ) ;
assign n1116 =  ( n1091 ) ? ( n387 ) : ( x21 ) ;
assign n1117 =  ( n1091 ) ? ( n393 ) : ( x21 ) ;
assign n1118 =  ( n1091 ) ? ( n395 ) : ( x21 ) ;
assign n1119 =  ( n230 ) ? ( n1118 ) : ( x21 ) ;
assign n1120 =  ( n229 ) ? ( n1117 ) : ( n1119 ) ;
assign n1121 =  ( n228 ) ? ( n1116 ) : ( n1120 ) ;
assign n1122 =  ( n227 ) ? ( n1115 ) : ( n1121 ) ;
assign n1123 =  ( n226 ) ? ( n1114 ) : ( n1122 ) ;
assign n1124 =  ( n220 ) ? ( n1113 ) : ( n1123 ) ;
assign n1125 =  ( n219 ) ? ( n1112 ) : ( n1124 ) ;
assign n1126 =  ( n343 ) ? ( n1111 ) : ( n1125 ) ;
assign n1127 =  ( n218 ) ? ( n1110 ) : ( n1126 ) ;
assign n1128 =  ( n217 ) ? ( n1109 ) : ( n1127 ) ;
assign n1129 =  ( n216 ) ? ( n1108 ) : ( n1128 ) ;
assign n1130 =  ( n215 ) ? ( n1107 ) : ( n1129 ) ;
assign n1131 =  ( n214 ) ? ( n1106 ) : ( n1130 ) ;
assign n1132 =  ( n213 ) ? ( n1105 ) : ( n1131 ) ;
assign n1133 =  ( n212 ) ? ( n1104 ) : ( n1132 ) ;
assign n1134 =  ( n210 ) ? ( n1103 ) : ( n1133 ) ;
assign n1135 =  ( n209 ) ? ( n1102 ) : ( n1134 ) ;
assign n1136 =  ( n206 ) ? ( n1101 ) : ( n1135 ) ;
assign n1137 =  ( n205 ) ? ( n1100 ) : ( n1136 ) ;
assign n1138 =  ( n202 ) ? ( n1099 ) : ( n1137 ) ;
assign n1139 =  ( n199 ) ? ( n1098 ) : ( n1138 ) ;
assign n1140 =  ( n197 ) ? ( n1097 ) : ( n1139 ) ;
assign n1141 =  ( n195 ) ? ( n1096 ) : ( n1140 ) ;
assign n1142 =  ( n193 ) ? ( n1095 ) : ( n1141 ) ;
assign n1143 =  ( n191 ) ? ( n1094 ) : ( n1142 ) ;
assign n1144 =  ( n189 ) ? ( n1093 ) : ( n1143 ) ;
assign n1145 =  ( n187 ) ? ( n1092 ) : ( n1144 ) ;
assign n1146 =  ( n296 ) == ( 5'd22 )  ;
assign n1147 =  ( n1146 ) ? ( n300 ) : ( x22 ) ;
assign n1148 =  ( n1146 ) ? ( n302 ) : ( x22 ) ;
assign n1149 =  ( n1146 ) ? ( n304 ) : ( x22 ) ;
assign n1150 =  ( n1146 ) ? ( n306 ) : ( x22 ) ;
assign n1151 =  ( n1146 ) ? ( n308 ) : ( x22 ) ;
assign n1152 =  ( n1146 ) ? ( n310 ) : ( x22 ) ;
assign n1153 =  ( n1146 ) ? ( n312 ) : ( x22 ) ;
assign n1154 =  ( n1146 ) ? ( n314 ) : ( x22 ) ;
assign n1155 =  ( n1146 ) ? ( n316 ) : ( x22 ) ;
assign n1156 =  ( n1146 ) ? ( n318 ) : ( x22 ) ;
assign n1157 =  ( n1146 ) ? ( n321 ) : ( x22 ) ;
assign n1158 =  ( n1146 ) ? ( n323 ) : ( x22 ) ;
assign n1159 =  ( n1146 ) ? ( n325 ) : ( x22 ) ;
assign n1160 =  ( n1146 ) ? ( n719 ) : ( x22 ) ;
assign n1161 =  ( n1146 ) ? ( n439 ) : ( x22 ) ;
assign n1162 =  ( n1146 ) ? ( n333 ) : ( x22 ) ;
assign n1163 =  ( n1146 ) ? ( n336 ) : ( x22 ) ;
assign n1164 =  ( n1146 ) ? ( n612 ) : ( x22 ) ;
assign n1165 =  ( n1146 ) ? ( n341 ) : ( x22 ) ;
assign n1166 =  ( n1146 ) ? ( n162 ) : ( x22 ) ;
assign n1167 =  ( n1146 ) ? ( n347 ) : ( x22 ) ;
assign n1168 =  ( n1146 ) ? ( n346 ) : ( x22 ) ;
assign n1169 =  ( n1146 ) ? ( n370 ) : ( x22 ) ;
assign n1170 =  ( n1146 ) ? ( n378 ) : ( x22 ) ;
assign n1171 =  ( n1146 ) ? ( n387 ) : ( x22 ) ;
assign n1172 =  ( n1146 ) ? ( n393 ) : ( x22 ) ;
assign n1173 =  ( n1146 ) ? ( n395 ) : ( x22 ) ;
assign n1174 =  ( n230 ) ? ( n1173 ) : ( x22 ) ;
assign n1175 =  ( n229 ) ? ( n1172 ) : ( n1174 ) ;
assign n1176 =  ( n228 ) ? ( n1171 ) : ( n1175 ) ;
assign n1177 =  ( n227 ) ? ( n1170 ) : ( n1176 ) ;
assign n1178 =  ( n226 ) ? ( n1169 ) : ( n1177 ) ;
assign n1179 =  ( n220 ) ? ( n1168 ) : ( n1178 ) ;
assign n1180 =  ( n219 ) ? ( n1167 ) : ( n1179 ) ;
assign n1181 =  ( n343 ) ? ( n1166 ) : ( n1180 ) ;
assign n1182 =  ( n218 ) ? ( n1165 ) : ( n1181 ) ;
assign n1183 =  ( n217 ) ? ( n1164 ) : ( n1182 ) ;
assign n1184 =  ( n216 ) ? ( n1163 ) : ( n1183 ) ;
assign n1185 =  ( n215 ) ? ( n1162 ) : ( n1184 ) ;
assign n1186 =  ( n214 ) ? ( n1161 ) : ( n1185 ) ;
assign n1187 =  ( n213 ) ? ( n1160 ) : ( n1186 ) ;
assign n1188 =  ( n212 ) ? ( n1159 ) : ( n1187 ) ;
assign n1189 =  ( n210 ) ? ( n1158 ) : ( n1188 ) ;
assign n1190 =  ( n209 ) ? ( n1157 ) : ( n1189 ) ;
assign n1191 =  ( n206 ) ? ( n1156 ) : ( n1190 ) ;
assign n1192 =  ( n205 ) ? ( n1155 ) : ( n1191 ) ;
assign n1193 =  ( n202 ) ? ( n1154 ) : ( n1192 ) ;
assign n1194 =  ( n199 ) ? ( n1153 ) : ( n1193 ) ;
assign n1195 =  ( n197 ) ? ( n1152 ) : ( n1194 ) ;
assign n1196 =  ( n195 ) ? ( n1151 ) : ( n1195 ) ;
assign n1197 =  ( n193 ) ? ( n1150 ) : ( n1196 ) ;
assign n1198 =  ( n191 ) ? ( n1149 ) : ( n1197 ) ;
assign n1199 =  ( n189 ) ? ( n1148 ) : ( n1198 ) ;
assign n1200 =  ( n187 ) ? ( n1147 ) : ( n1199 ) ;
assign n1201 =  ( n296 ) == ( 5'd23 )  ;
assign n1202 =  ( n1201 ) ? ( n300 ) : ( x23 ) ;
assign n1203 =  ( n1201 ) ? ( n302 ) : ( x23 ) ;
assign n1204 =  ( n1201 ) ? ( n304 ) : ( x23 ) ;
assign n1205 =  ( n1201 ) ? ( n306 ) : ( x23 ) ;
assign n1206 =  ( n1201 ) ? ( n308 ) : ( x23 ) ;
assign n1207 =  ( n1201 ) ? ( n310 ) : ( x23 ) ;
assign n1208 =  ( n1201 ) ? ( n312 ) : ( x23 ) ;
assign n1209 =  ( n1201 ) ? ( n314 ) : ( x23 ) ;
assign n1210 =  ( n1201 ) ? ( n316 ) : ( x23 ) ;
assign n1211 =  ( n1201 ) ? ( n318 ) : ( x23 ) ;
assign n1212 =  ( n1201 ) ? ( n321 ) : ( x23 ) ;
assign n1213 =  ( n1201 ) ? ( n323 ) : ( x23 ) ;
assign n1214 =  ( n1201 ) ? ( n325 ) : ( x23 ) ;
assign n1215 =  ( n1201 ) ? ( n719 ) : ( x23 ) ;
assign n1216 =  ( n1201 ) ? ( n439 ) : ( x23 ) ;
assign n1217 =  ( n1201 ) ? ( n333 ) : ( x23 ) ;
assign n1218 =  ( n1201 ) ? ( n553 ) : ( x23 ) ;
assign n1219 =  ( n1201 ) ? ( n612 ) : ( x23 ) ;
assign n1220 =  ( n1201 ) ? ( n341 ) : ( x23 ) ;
assign n1221 =  ( n1201 ) ? ( n162 ) : ( x23 ) ;
assign n1222 =  ( n1201 ) ? ( n347 ) : ( x23 ) ;
assign n1223 =  ( n1201 ) ? ( n346 ) : ( x23 ) ;
assign n1224 =  ( n1201 ) ? ( n370 ) : ( x23 ) ;
assign n1225 =  ( n1201 ) ? ( n378 ) : ( x23 ) ;
assign n1226 =  ( n1201 ) ? ( n387 ) : ( x23 ) ;
assign n1227 =  ( n1201 ) ? ( n393 ) : ( x23 ) ;
assign n1228 =  ( n1201 ) ? ( n395 ) : ( x23 ) ;
assign n1229 =  ( n230 ) ? ( n1228 ) : ( x23 ) ;
assign n1230 =  ( n229 ) ? ( n1227 ) : ( n1229 ) ;
assign n1231 =  ( n228 ) ? ( n1226 ) : ( n1230 ) ;
assign n1232 =  ( n227 ) ? ( n1225 ) : ( n1231 ) ;
assign n1233 =  ( n226 ) ? ( n1224 ) : ( n1232 ) ;
assign n1234 =  ( n220 ) ? ( n1223 ) : ( n1233 ) ;
assign n1235 =  ( n219 ) ? ( n1222 ) : ( n1234 ) ;
assign n1236 =  ( n343 ) ? ( n1221 ) : ( n1235 ) ;
assign n1237 =  ( n218 ) ? ( n1220 ) : ( n1236 ) ;
assign n1238 =  ( n217 ) ? ( n1219 ) : ( n1237 ) ;
assign n1239 =  ( n216 ) ? ( n1218 ) : ( n1238 ) ;
assign n1240 =  ( n215 ) ? ( n1217 ) : ( n1239 ) ;
assign n1241 =  ( n214 ) ? ( n1216 ) : ( n1240 ) ;
assign n1242 =  ( n213 ) ? ( n1215 ) : ( n1241 ) ;
assign n1243 =  ( n212 ) ? ( n1214 ) : ( n1242 ) ;
assign n1244 =  ( n210 ) ? ( n1213 ) : ( n1243 ) ;
assign n1245 =  ( n209 ) ? ( n1212 ) : ( n1244 ) ;
assign n1246 =  ( n206 ) ? ( n1211 ) : ( n1245 ) ;
assign n1247 =  ( n205 ) ? ( n1210 ) : ( n1246 ) ;
assign n1248 =  ( n202 ) ? ( n1209 ) : ( n1247 ) ;
assign n1249 =  ( n199 ) ? ( n1208 ) : ( n1248 ) ;
assign n1250 =  ( n197 ) ? ( n1207 ) : ( n1249 ) ;
assign n1251 =  ( n195 ) ? ( n1206 ) : ( n1250 ) ;
assign n1252 =  ( n193 ) ? ( n1205 ) : ( n1251 ) ;
assign n1253 =  ( n191 ) ? ( n1204 ) : ( n1252 ) ;
assign n1254 =  ( n189 ) ? ( n1203 ) : ( n1253 ) ;
assign n1255 =  ( n187 ) ? ( n1202 ) : ( n1254 ) ;
assign n1256 =  ( n296 ) == ( 5'd24 )  ;
assign n1257 =  ( n1256 ) ? ( n300 ) : ( x24 ) ;
assign n1258 =  ( n1256 ) ? ( n302 ) : ( x24 ) ;
assign n1259 =  ( n1256 ) ? ( n304 ) : ( x24 ) ;
assign n1260 =  ( n1256 ) ? ( n306 ) : ( x24 ) ;
assign n1261 =  ( n1256 ) ? ( n308 ) : ( x24 ) ;
assign n1262 =  ( n1256 ) ? ( n310 ) : ( x24 ) ;
assign n1263 =  ( n1256 ) ? ( n312 ) : ( x24 ) ;
assign n1264 =  ( n1256 ) ? ( n314 ) : ( x24 ) ;
assign n1265 =  ( n1256 ) ? ( n316 ) : ( x24 ) ;
assign n1266 =  ( n1256 ) ? ( n318 ) : ( x24 ) ;
assign n1267 =  ( n1256 ) ? ( n321 ) : ( x24 ) ;
assign n1268 =  ( n1256 ) ? ( n323 ) : ( x24 ) ;
assign n1269 =  ( n1256 ) ? ( n325 ) : ( x24 ) ;
assign n1270 =  ( n1256 ) ? ( n328 ) : ( x24 ) ;
assign n1271 =  ( n1256 ) ? ( n439 ) : ( x24 ) ;
assign n1272 =  ( n1256 ) ? ( n333 ) : ( x24 ) ;
assign n1273 =  ( n1256 ) ? ( n553 ) : ( x24 ) ;
assign n1274 =  ( n1256 ) ? ( n339 ) : ( x24 ) ;
assign n1275 =  ( n1256 ) ? ( n341 ) : ( x24 ) ;
assign n1276 =  ( n1256 ) ? ( n162 ) : ( x24 ) ;
assign n1277 =  ( n1256 ) ? ( n347 ) : ( x24 ) ;
assign n1278 =  ( n1256 ) ? ( n346 ) : ( x24 ) ;
assign n1279 =  ( n1256 ) ? ( n370 ) : ( x24 ) ;
assign n1280 =  ( n1256 ) ? ( n378 ) : ( x24 ) ;
assign n1281 =  ( n1256 ) ? ( n387 ) : ( x24 ) ;
assign n1282 =  ( n1256 ) ? ( n393 ) : ( x24 ) ;
assign n1283 =  ( n1256 ) ? ( n395 ) : ( x24 ) ;
assign n1284 =  ( n230 ) ? ( n1283 ) : ( x24 ) ;
assign n1285 =  ( n229 ) ? ( n1282 ) : ( n1284 ) ;
assign n1286 =  ( n228 ) ? ( n1281 ) : ( n1285 ) ;
assign n1287 =  ( n227 ) ? ( n1280 ) : ( n1286 ) ;
assign n1288 =  ( n226 ) ? ( n1279 ) : ( n1287 ) ;
assign n1289 =  ( n220 ) ? ( n1278 ) : ( n1288 ) ;
assign n1290 =  ( n219 ) ? ( n1277 ) : ( n1289 ) ;
assign n1291 =  ( n343 ) ? ( n1276 ) : ( n1290 ) ;
assign n1292 =  ( n218 ) ? ( n1275 ) : ( n1291 ) ;
assign n1293 =  ( n217 ) ? ( n1274 ) : ( n1292 ) ;
assign n1294 =  ( n216 ) ? ( n1273 ) : ( n1293 ) ;
assign n1295 =  ( n215 ) ? ( n1272 ) : ( n1294 ) ;
assign n1296 =  ( n214 ) ? ( n1271 ) : ( n1295 ) ;
assign n1297 =  ( n213 ) ? ( n1270 ) : ( n1296 ) ;
assign n1298 =  ( n212 ) ? ( n1269 ) : ( n1297 ) ;
assign n1299 =  ( n210 ) ? ( n1268 ) : ( n1298 ) ;
assign n1300 =  ( n209 ) ? ( n1267 ) : ( n1299 ) ;
assign n1301 =  ( n206 ) ? ( n1266 ) : ( n1300 ) ;
assign n1302 =  ( n205 ) ? ( n1265 ) : ( n1301 ) ;
assign n1303 =  ( n202 ) ? ( n1264 ) : ( n1302 ) ;
assign n1304 =  ( n199 ) ? ( n1263 ) : ( n1303 ) ;
assign n1305 =  ( n197 ) ? ( n1262 ) : ( n1304 ) ;
assign n1306 =  ( n195 ) ? ( n1261 ) : ( n1305 ) ;
assign n1307 =  ( n193 ) ? ( n1260 ) : ( n1306 ) ;
assign n1308 =  ( n191 ) ? ( n1259 ) : ( n1307 ) ;
assign n1309 =  ( n189 ) ? ( n1258 ) : ( n1308 ) ;
assign n1310 =  ( n187 ) ? ( n1257 ) : ( n1309 ) ;
assign n1311 =  ( n296 ) == ( 5'd25 )  ;
assign n1312 =  ( n1311 ) ? ( n300 ) : ( x25 ) ;
assign n1313 =  ( n1311 ) ? ( n302 ) : ( x25 ) ;
assign n1314 =  ( n1311 ) ? ( n304 ) : ( x25 ) ;
assign n1315 =  ( n1311 ) ? ( n306 ) : ( x25 ) ;
assign n1316 =  ( n1311 ) ? ( n308 ) : ( x25 ) ;
assign n1317 =  ( n1311 ) ? ( n310 ) : ( x25 ) ;
assign n1318 =  ( n1311 ) ? ( n312 ) : ( x25 ) ;
assign n1319 =  ( n1311 ) ? ( n314 ) : ( x25 ) ;
assign n1320 =  ( n1311 ) ? ( n316 ) : ( x25 ) ;
assign n1321 =  ( n1311 ) ? ( n318 ) : ( x25 ) ;
assign n1322 =  ( n1311 ) ? ( n321 ) : ( x25 ) ;
assign n1323 =  ( n1311 ) ? ( n323 ) : ( x25 ) ;
assign n1324 =  ( n1311 ) ? ( n325 ) : ( x25 ) ;
assign n1325 =  ( n1311 ) ? ( n328 ) : ( x25 ) ;
assign n1326 =  ( n1311 ) ? ( n439 ) : ( x25 ) ;
assign n1327 =  ( n1311 ) ? ( n333 ) : ( x25 ) ;
assign n1328 =  ( n1311 ) ? ( n336 ) : ( x25 ) ;
assign n1329 =  ( n1311 ) ? ( n339 ) : ( x25 ) ;
assign n1330 =  ( n1311 ) ? ( n341 ) : ( x25 ) ;
assign n1331 =  ( n1311 ) ? ( n162 ) : ( x25 ) ;
assign n1332 =  ( n1311 ) ? ( n347 ) : ( x25 ) ;
assign n1333 =  ( n1311 ) ? ( n346 ) : ( x25 ) ;
assign n1334 =  ( n1311 ) ? ( n370 ) : ( x25 ) ;
assign n1335 =  ( n1311 ) ? ( n378 ) : ( x25 ) ;
assign n1336 =  ( n1311 ) ? ( n387 ) : ( x25 ) ;
assign n1337 =  ( n1311 ) ? ( n393 ) : ( x25 ) ;
assign n1338 =  ( n1311 ) ? ( n395 ) : ( x25 ) ;
assign n1339 =  ( n230 ) ? ( n1338 ) : ( x25 ) ;
assign n1340 =  ( n229 ) ? ( n1337 ) : ( n1339 ) ;
assign n1341 =  ( n228 ) ? ( n1336 ) : ( n1340 ) ;
assign n1342 =  ( n227 ) ? ( n1335 ) : ( n1341 ) ;
assign n1343 =  ( n226 ) ? ( n1334 ) : ( n1342 ) ;
assign n1344 =  ( n220 ) ? ( n1333 ) : ( n1343 ) ;
assign n1345 =  ( n219 ) ? ( n1332 ) : ( n1344 ) ;
assign n1346 =  ( n343 ) ? ( n1331 ) : ( n1345 ) ;
assign n1347 =  ( n218 ) ? ( n1330 ) : ( n1346 ) ;
assign n1348 =  ( n217 ) ? ( n1329 ) : ( n1347 ) ;
assign n1349 =  ( n216 ) ? ( n1328 ) : ( n1348 ) ;
assign n1350 =  ( n215 ) ? ( n1327 ) : ( n1349 ) ;
assign n1351 =  ( n214 ) ? ( n1326 ) : ( n1350 ) ;
assign n1352 =  ( n213 ) ? ( n1325 ) : ( n1351 ) ;
assign n1353 =  ( n212 ) ? ( n1324 ) : ( n1352 ) ;
assign n1354 =  ( n210 ) ? ( n1323 ) : ( n1353 ) ;
assign n1355 =  ( n209 ) ? ( n1322 ) : ( n1354 ) ;
assign n1356 =  ( n206 ) ? ( n1321 ) : ( n1355 ) ;
assign n1357 =  ( n205 ) ? ( n1320 ) : ( n1356 ) ;
assign n1358 =  ( n202 ) ? ( n1319 ) : ( n1357 ) ;
assign n1359 =  ( n199 ) ? ( n1318 ) : ( n1358 ) ;
assign n1360 =  ( n197 ) ? ( n1317 ) : ( n1359 ) ;
assign n1361 =  ( n195 ) ? ( n1316 ) : ( n1360 ) ;
assign n1362 =  ( n193 ) ? ( n1315 ) : ( n1361 ) ;
assign n1363 =  ( n191 ) ? ( n1314 ) : ( n1362 ) ;
assign n1364 =  ( n189 ) ? ( n1313 ) : ( n1363 ) ;
assign n1365 =  ( n187 ) ? ( n1312 ) : ( n1364 ) ;
assign n1366 =  ( n296 ) == ( 5'd26 )  ;
assign n1367 =  ( n1366 ) ? ( n300 ) : ( x26 ) ;
assign n1368 =  ( n1366 ) ? ( n302 ) : ( x26 ) ;
assign n1369 =  ( n1366 ) ? ( n304 ) : ( x26 ) ;
assign n1370 =  ( n1366 ) ? ( n306 ) : ( x26 ) ;
assign n1371 =  ( n1366 ) ? ( n308 ) : ( x26 ) ;
assign n1372 =  ( n1366 ) ? ( n310 ) : ( x26 ) ;
assign n1373 =  ( n1366 ) ? ( n312 ) : ( x26 ) ;
assign n1374 =  ( n1366 ) ? ( n314 ) : ( x26 ) ;
assign n1375 =  ( n1366 ) ? ( n316 ) : ( x26 ) ;
assign n1376 =  ( n1366 ) ? ( n318 ) : ( x26 ) ;
assign n1377 =  ( n1366 ) ? ( n321 ) : ( x26 ) ;
assign n1378 =  ( n1366 ) ? ( n323 ) : ( x26 ) ;
assign n1379 =  ( n1366 ) ? ( n325 ) : ( x26 ) ;
assign n1380 =  ( n1366 ) ? ( n328 ) : ( x26 ) ;
assign n1381 =  ( n1366 ) ? ( n439 ) : ( x26 ) ;
assign n1382 =  ( n1366 ) ? ( n333 ) : ( x26 ) ;
assign n1383 =  ( n1366 ) ? ( n553 ) : ( x26 ) ;
assign n1384 =  ( n1366 ) ? ( n339 ) : ( x26 ) ;
assign n1385 =  ( n1366 ) ? ( n341 ) : ( x26 ) ;
assign n1386 =  ( n1366 ) ? ( n162 ) : ( x26 ) ;
assign n1387 =  ( n1366 ) ? ( n347 ) : ( x26 ) ;
assign n1388 =  ( n1366 ) ? ( n346 ) : ( x26 ) ;
assign n1389 =  ( n1366 ) ? ( n370 ) : ( x26 ) ;
assign n1390 =  ( n1366 ) ? ( n378 ) : ( x26 ) ;
assign n1391 =  ( n1366 ) ? ( n387 ) : ( x26 ) ;
assign n1392 =  ( n1366 ) ? ( n393 ) : ( x26 ) ;
assign n1393 =  ( n1366 ) ? ( n395 ) : ( x26 ) ;
assign n1394 =  ( n230 ) ? ( n1393 ) : ( x26 ) ;
assign n1395 =  ( n229 ) ? ( n1392 ) : ( n1394 ) ;
assign n1396 =  ( n228 ) ? ( n1391 ) : ( n1395 ) ;
assign n1397 =  ( n227 ) ? ( n1390 ) : ( n1396 ) ;
assign n1398 =  ( n226 ) ? ( n1389 ) : ( n1397 ) ;
assign n1399 =  ( n220 ) ? ( n1388 ) : ( n1398 ) ;
assign n1400 =  ( n219 ) ? ( n1387 ) : ( n1399 ) ;
assign n1401 =  ( n343 ) ? ( n1386 ) : ( n1400 ) ;
assign n1402 =  ( n218 ) ? ( n1385 ) : ( n1401 ) ;
assign n1403 =  ( n217 ) ? ( n1384 ) : ( n1402 ) ;
assign n1404 =  ( n216 ) ? ( n1383 ) : ( n1403 ) ;
assign n1405 =  ( n215 ) ? ( n1382 ) : ( n1404 ) ;
assign n1406 =  ( n214 ) ? ( n1381 ) : ( n1405 ) ;
assign n1407 =  ( n213 ) ? ( n1380 ) : ( n1406 ) ;
assign n1408 =  ( n212 ) ? ( n1379 ) : ( n1407 ) ;
assign n1409 =  ( n210 ) ? ( n1378 ) : ( n1408 ) ;
assign n1410 =  ( n209 ) ? ( n1377 ) : ( n1409 ) ;
assign n1411 =  ( n206 ) ? ( n1376 ) : ( n1410 ) ;
assign n1412 =  ( n205 ) ? ( n1375 ) : ( n1411 ) ;
assign n1413 =  ( n202 ) ? ( n1374 ) : ( n1412 ) ;
assign n1414 =  ( n199 ) ? ( n1373 ) : ( n1413 ) ;
assign n1415 =  ( n197 ) ? ( n1372 ) : ( n1414 ) ;
assign n1416 =  ( n195 ) ? ( n1371 ) : ( n1415 ) ;
assign n1417 =  ( n193 ) ? ( n1370 ) : ( n1416 ) ;
assign n1418 =  ( n191 ) ? ( n1369 ) : ( n1417 ) ;
assign n1419 =  ( n189 ) ? ( n1368 ) : ( n1418 ) ;
assign n1420 =  ( n187 ) ? ( n1367 ) : ( n1419 ) ;
assign n1421 =  ( n296 ) == ( 5'd27 )  ;
assign n1422 =  ( n1421 ) ? ( n300 ) : ( x27 ) ;
assign n1423 =  ( n1421 ) ? ( n302 ) : ( x27 ) ;
assign n1424 =  ( n1421 ) ? ( n304 ) : ( x27 ) ;
assign n1425 =  ( n1421 ) ? ( n306 ) : ( x27 ) ;
assign n1426 =  ( n1421 ) ? ( n308 ) : ( x27 ) ;
assign n1427 =  ( n1421 ) ? ( n310 ) : ( x27 ) ;
assign n1428 =  ( n1421 ) ? ( n312 ) : ( x27 ) ;
assign n1429 =  ( n1421 ) ? ( n314 ) : ( x27 ) ;
assign n1430 =  ( n1421 ) ? ( n316 ) : ( x27 ) ;
assign n1431 =  ( n1421 ) ? ( n318 ) : ( x27 ) ;
assign n1432 =  ( n1421 ) ? ( n321 ) : ( x27 ) ;
assign n1433 =  ( n1421 ) ? ( n323 ) : ( x27 ) ;
assign n1434 =  ( n1421 ) ? ( n325 ) : ( x27 ) ;
assign n1435 =  ( n1421 ) ? ( n328 ) : ( x27 ) ;
assign n1436 =  ( n1421 ) ? ( n439 ) : ( x27 ) ;
assign n1437 =  ( n1421 ) ? ( n608 ) : ( x27 ) ;
assign n1438 =  ( n1421 ) ? ( n336 ) : ( x27 ) ;
assign n1439 =  ( n1421 ) ? ( n339 ) : ( x27 ) ;
assign n1440 =  ( n1421 ) ? ( n341 ) : ( x27 ) ;
assign n1441 =  ( n1421 ) ? ( n162 ) : ( x27 ) ;
assign n1442 =  ( n1421 ) ? ( n347 ) : ( x27 ) ;
assign n1443 =  ( n1421 ) ? ( n346 ) : ( x27 ) ;
assign n1444 =  ( n1421 ) ? ( n370 ) : ( x27 ) ;
assign n1445 =  ( n1421 ) ? ( n378 ) : ( x27 ) ;
assign n1446 =  ( n1421 ) ? ( n387 ) : ( x27 ) ;
assign n1447 =  ( n1421 ) ? ( n393 ) : ( x27 ) ;
assign n1448 =  ( n1421 ) ? ( n395 ) : ( x27 ) ;
assign n1449 =  ( n230 ) ? ( n1448 ) : ( x27 ) ;
assign n1450 =  ( n229 ) ? ( n1447 ) : ( n1449 ) ;
assign n1451 =  ( n228 ) ? ( n1446 ) : ( n1450 ) ;
assign n1452 =  ( n227 ) ? ( n1445 ) : ( n1451 ) ;
assign n1453 =  ( n226 ) ? ( n1444 ) : ( n1452 ) ;
assign n1454 =  ( n220 ) ? ( n1443 ) : ( n1453 ) ;
assign n1455 =  ( n219 ) ? ( n1442 ) : ( n1454 ) ;
assign n1456 =  ( n343 ) ? ( n1441 ) : ( n1455 ) ;
assign n1457 =  ( n218 ) ? ( n1440 ) : ( n1456 ) ;
assign n1458 =  ( n217 ) ? ( n1439 ) : ( n1457 ) ;
assign n1459 =  ( n216 ) ? ( n1438 ) : ( n1458 ) ;
assign n1460 =  ( n215 ) ? ( n1437 ) : ( n1459 ) ;
assign n1461 =  ( n214 ) ? ( n1436 ) : ( n1460 ) ;
assign n1462 =  ( n213 ) ? ( n1435 ) : ( n1461 ) ;
assign n1463 =  ( n212 ) ? ( n1434 ) : ( n1462 ) ;
assign n1464 =  ( n210 ) ? ( n1433 ) : ( n1463 ) ;
assign n1465 =  ( n209 ) ? ( n1432 ) : ( n1464 ) ;
assign n1466 =  ( n206 ) ? ( n1431 ) : ( n1465 ) ;
assign n1467 =  ( n205 ) ? ( n1430 ) : ( n1466 ) ;
assign n1468 =  ( n202 ) ? ( n1429 ) : ( n1467 ) ;
assign n1469 =  ( n199 ) ? ( n1428 ) : ( n1468 ) ;
assign n1470 =  ( n197 ) ? ( n1427 ) : ( n1469 ) ;
assign n1471 =  ( n195 ) ? ( n1426 ) : ( n1470 ) ;
assign n1472 =  ( n193 ) ? ( n1425 ) : ( n1471 ) ;
assign n1473 =  ( n191 ) ? ( n1424 ) : ( n1472 ) ;
assign n1474 =  ( n189 ) ? ( n1423 ) : ( n1473 ) ;
assign n1475 =  ( n187 ) ? ( n1422 ) : ( n1474 ) ;
assign n1476 =  ( n296 ) == ( 5'd28 )  ;
assign n1477 =  ( n1476 ) ? ( n300 ) : ( x28 ) ;
assign n1478 =  ( n1476 ) ? ( n302 ) : ( x28 ) ;
assign n1479 =  ( n1476 ) ? ( n304 ) : ( x28 ) ;
assign n1480 =  ( n1476 ) ? ( n306 ) : ( x28 ) ;
assign n1481 =  ( n1476 ) ? ( n308 ) : ( x28 ) ;
assign n1482 =  ( n1476 ) ? ( n310 ) : ( x28 ) ;
assign n1483 =  ( n1476 ) ? ( n312 ) : ( x28 ) ;
assign n1484 =  ( n1476 ) ? ( n314 ) : ( x28 ) ;
assign n1485 =  ( n1476 ) ? ( n316 ) : ( x28 ) ;
assign n1486 =  ( n1476 ) ? ( n318 ) : ( x28 ) ;
assign n1487 =  ( n1476 ) ? ( n321 ) : ( x28 ) ;
assign n1488 =  ( n1476 ) ? ( n323 ) : ( x28 ) ;
assign n1489 =  ( n1476 ) ? ( n325 ) : ( x28 ) ;
assign n1490 =  ( n1476 ) ? ( n328 ) : ( x28 ) ;
assign n1491 =  ( n1476 ) ? ( n439 ) : ( x28 ) ;
assign n1492 =  ( n1476 ) ? ( n333 ) : ( x28 ) ;
assign n1493 =  ( n1476 ) ? ( n336 ) : ( x28 ) ;
assign n1494 =  ( n1476 ) ? ( n339 ) : ( x28 ) ;
assign n1495 =  ( n1476 ) ? ( n341 ) : ( x28 ) ;
assign n1496 =  ( n1476 ) ? ( n162 ) : ( x28 ) ;
assign n1497 =  ( n1476 ) ? ( n347 ) : ( x28 ) ;
assign n1498 =  ( n1476 ) ? ( n346 ) : ( x28 ) ;
assign n1499 =  ( n1476 ) ? ( n370 ) : ( x28 ) ;
assign n1500 =  ( n1476 ) ? ( n378 ) : ( x28 ) ;
assign n1501 =  ( n1476 ) ? ( n387 ) : ( x28 ) ;
assign n1502 =  ( n1476 ) ? ( n393 ) : ( x28 ) ;
assign n1503 =  ( n1476 ) ? ( n395 ) : ( x28 ) ;
assign n1504 =  ( n230 ) ? ( n1503 ) : ( x28 ) ;
assign n1505 =  ( n229 ) ? ( n1502 ) : ( n1504 ) ;
assign n1506 =  ( n228 ) ? ( n1501 ) : ( n1505 ) ;
assign n1507 =  ( n227 ) ? ( n1500 ) : ( n1506 ) ;
assign n1508 =  ( n226 ) ? ( n1499 ) : ( n1507 ) ;
assign n1509 =  ( n220 ) ? ( n1498 ) : ( n1508 ) ;
assign n1510 =  ( n219 ) ? ( n1497 ) : ( n1509 ) ;
assign n1511 =  ( n343 ) ? ( n1496 ) : ( n1510 ) ;
assign n1512 =  ( n218 ) ? ( n1495 ) : ( n1511 ) ;
assign n1513 =  ( n217 ) ? ( n1494 ) : ( n1512 ) ;
assign n1514 =  ( n216 ) ? ( n1493 ) : ( n1513 ) ;
assign n1515 =  ( n215 ) ? ( n1492 ) : ( n1514 ) ;
assign n1516 =  ( n214 ) ? ( n1491 ) : ( n1515 ) ;
assign n1517 =  ( n213 ) ? ( n1490 ) : ( n1516 ) ;
assign n1518 =  ( n212 ) ? ( n1489 ) : ( n1517 ) ;
assign n1519 =  ( n210 ) ? ( n1488 ) : ( n1518 ) ;
assign n1520 =  ( n209 ) ? ( n1487 ) : ( n1519 ) ;
assign n1521 =  ( n206 ) ? ( n1486 ) : ( n1520 ) ;
assign n1522 =  ( n205 ) ? ( n1485 ) : ( n1521 ) ;
assign n1523 =  ( n202 ) ? ( n1484 ) : ( n1522 ) ;
assign n1524 =  ( n199 ) ? ( n1483 ) : ( n1523 ) ;
assign n1525 =  ( n197 ) ? ( n1482 ) : ( n1524 ) ;
assign n1526 =  ( n195 ) ? ( n1481 ) : ( n1525 ) ;
assign n1527 =  ( n193 ) ? ( n1480 ) : ( n1526 ) ;
assign n1528 =  ( n191 ) ? ( n1479 ) : ( n1527 ) ;
assign n1529 =  ( n189 ) ? ( n1478 ) : ( n1528 ) ;
assign n1530 =  ( n187 ) ? ( n1477 ) : ( n1529 ) ;
assign n1531 =  ( n296 ) == ( 5'd29 )  ;
assign n1532 =  ( n1531 ) ? ( n300 ) : ( x29 ) ;
assign n1533 =  ( n1531 ) ? ( n302 ) : ( x29 ) ;
assign n1534 =  ( n1531 ) ? ( n304 ) : ( x29 ) ;
assign n1535 =  ( n1531 ) ? ( n306 ) : ( x29 ) ;
assign n1536 =  ( n1531 ) ? ( n308 ) : ( x29 ) ;
assign n1537 =  ( n1531 ) ? ( n310 ) : ( x29 ) ;
assign n1538 =  ( n1531 ) ? ( n312 ) : ( x29 ) ;
assign n1539 =  ( n1531 ) ? ( n314 ) : ( x29 ) ;
assign n1540 =  ( n1531 ) ? ( n316 ) : ( x29 ) ;
assign n1541 =  ( n1531 ) ? ( n318 ) : ( x29 ) ;
assign n1542 =  ( n1531 ) ? ( n321 ) : ( x29 ) ;
assign n1543 =  ( n1531 ) ? ( n323 ) : ( x29 ) ;
assign n1544 =  ( n1531 ) ? ( n325 ) : ( x29 ) ;
assign n1545 =  ( n1531 ) ? ( n328 ) : ( x29 ) ;
assign n1546 =  ( n1531 ) ? ( n439 ) : ( x29 ) ;
assign n1547 =  ( n1531 ) ? ( n608 ) : ( x29 ) ;
assign n1548 =  ( n1531 ) ? ( n553 ) : ( x29 ) ;
assign n1549 =  ( n1531 ) ? ( n612 ) : ( x29 ) ;
assign n1550 =  ( n1531 ) ? ( n341 ) : ( x29 ) ;
assign n1551 =  ( n1531 ) ? ( n162 ) : ( x29 ) ;
assign n1552 =  ( n1531 ) ? ( n347 ) : ( x29 ) ;
assign n1553 =  ( n1531 ) ? ( n346 ) : ( x29 ) ;
assign n1554 =  ( n1531 ) ? ( n370 ) : ( x29 ) ;
assign n1555 =  ( n1531 ) ? ( n378 ) : ( x29 ) ;
assign n1556 =  ( n1531 ) ? ( n387 ) : ( x29 ) ;
assign n1557 =  ( n1531 ) ? ( n393 ) : ( x29 ) ;
assign n1558 =  ( n1531 ) ? ( n395 ) : ( x29 ) ;
assign n1559 =  ( n230 ) ? ( n1558 ) : ( x29 ) ;
assign n1560 =  ( n229 ) ? ( n1557 ) : ( n1559 ) ;
assign n1561 =  ( n228 ) ? ( n1556 ) : ( n1560 ) ;
assign n1562 =  ( n227 ) ? ( n1555 ) : ( n1561 ) ;
assign n1563 =  ( n226 ) ? ( n1554 ) : ( n1562 ) ;
assign n1564 =  ( n220 ) ? ( n1553 ) : ( n1563 ) ;
assign n1565 =  ( n219 ) ? ( n1552 ) : ( n1564 ) ;
assign n1566 =  ( n343 ) ? ( n1551 ) : ( n1565 ) ;
assign n1567 =  ( n218 ) ? ( n1550 ) : ( n1566 ) ;
assign n1568 =  ( n217 ) ? ( n1549 ) : ( n1567 ) ;
assign n1569 =  ( n216 ) ? ( n1548 ) : ( n1568 ) ;
assign n1570 =  ( n215 ) ? ( n1547 ) : ( n1569 ) ;
assign n1571 =  ( n214 ) ? ( n1546 ) : ( n1570 ) ;
assign n1572 =  ( n213 ) ? ( n1545 ) : ( n1571 ) ;
assign n1573 =  ( n212 ) ? ( n1544 ) : ( n1572 ) ;
assign n1574 =  ( n210 ) ? ( n1543 ) : ( n1573 ) ;
assign n1575 =  ( n209 ) ? ( n1542 ) : ( n1574 ) ;
assign n1576 =  ( n206 ) ? ( n1541 ) : ( n1575 ) ;
assign n1577 =  ( n205 ) ? ( n1540 ) : ( n1576 ) ;
assign n1578 =  ( n202 ) ? ( n1539 ) : ( n1577 ) ;
assign n1579 =  ( n199 ) ? ( n1538 ) : ( n1578 ) ;
assign n1580 =  ( n197 ) ? ( n1537 ) : ( n1579 ) ;
assign n1581 =  ( n195 ) ? ( n1536 ) : ( n1580 ) ;
assign n1582 =  ( n193 ) ? ( n1535 ) : ( n1581 ) ;
assign n1583 =  ( n191 ) ? ( n1534 ) : ( n1582 ) ;
assign n1584 =  ( n189 ) ? ( n1533 ) : ( n1583 ) ;
assign n1585 =  ( n187 ) ? ( n1532 ) : ( n1584 ) ;
assign n1586 =  ( n296 ) == ( 5'd3 )  ;
assign n1587 =  ( n1586 ) ? ( n300 ) : ( x3 ) ;
assign n1588 =  ( n1586 ) ? ( n302 ) : ( x3 ) ;
assign n1589 =  ( n1586 ) ? ( n304 ) : ( x3 ) ;
assign n1590 =  ( n1586 ) ? ( n306 ) : ( x3 ) ;
assign n1591 =  ( n1586 ) ? ( n308 ) : ( x3 ) ;
assign n1592 =  ( n1586 ) ? ( n310 ) : ( x3 ) ;
assign n1593 =  ( n1586 ) ? ( n312 ) : ( x3 ) ;
assign n1594 =  ( n1586 ) ? ( n314 ) : ( x3 ) ;
assign n1595 =  ( n1586 ) ? ( n316 ) : ( x3 ) ;
assign n1596 =  ( n1586 ) ? ( n318 ) : ( x3 ) ;
assign n1597 =  ( n1586 ) ? ( n321 ) : ( x3 ) ;
assign n1598 =  ( n1586 ) ? ( n323 ) : ( x3 ) ;
assign n1599 =  ( n1586 ) ? ( n325 ) : ( x3 ) ;
assign n1600 =  ( n1586 ) ? ( n328 ) : ( x3 ) ;
assign n1601 =  ( n1586 ) ? ( n439 ) : ( x3 ) ;
assign n1602 =  ( n1586 ) ? ( n608 ) : ( x3 ) ;
assign n1603 =  ( n1586 ) ? ( n336 ) : ( x3 ) ;
assign n1604 =  ( n1586 ) ? ( n339 ) : ( x3 ) ;
assign n1605 =  ( n1586 ) ? ( n341 ) : ( x3 ) ;
assign n1606 =  ( n1586 ) ? ( n162 ) : ( x3 ) ;
assign n1607 =  ( n1586 ) ? ( n347 ) : ( x3 ) ;
assign n1608 =  ( n1586 ) ? ( n346 ) : ( x3 ) ;
assign n1609 =  ( n1586 ) ? ( n370 ) : ( x3 ) ;
assign n1610 =  ( n1586 ) ? ( n378 ) : ( x3 ) ;
assign n1611 =  ( n1586 ) ? ( n387 ) : ( x3 ) ;
assign n1612 =  ( n1586 ) ? ( n393 ) : ( x3 ) ;
assign n1613 =  ( n1586 ) ? ( n395 ) : ( x3 ) ;
assign n1614 =  ( n230 ) ? ( n1613 ) : ( x3 ) ;
assign n1615 =  ( n229 ) ? ( n1612 ) : ( n1614 ) ;
assign n1616 =  ( n228 ) ? ( n1611 ) : ( n1615 ) ;
assign n1617 =  ( n227 ) ? ( n1610 ) : ( n1616 ) ;
assign n1618 =  ( n226 ) ? ( n1609 ) : ( n1617 ) ;
assign n1619 =  ( n220 ) ? ( n1608 ) : ( n1618 ) ;
assign n1620 =  ( n219 ) ? ( n1607 ) : ( n1619 ) ;
assign n1621 =  ( n343 ) ? ( n1606 ) : ( n1620 ) ;
assign n1622 =  ( n218 ) ? ( n1605 ) : ( n1621 ) ;
assign n1623 =  ( n217 ) ? ( n1604 ) : ( n1622 ) ;
assign n1624 =  ( n216 ) ? ( n1603 ) : ( n1623 ) ;
assign n1625 =  ( n215 ) ? ( n1602 ) : ( n1624 ) ;
assign n1626 =  ( n214 ) ? ( n1601 ) : ( n1625 ) ;
assign n1627 =  ( n213 ) ? ( n1600 ) : ( n1626 ) ;
assign n1628 =  ( n212 ) ? ( n1599 ) : ( n1627 ) ;
assign n1629 =  ( n210 ) ? ( n1598 ) : ( n1628 ) ;
assign n1630 =  ( n209 ) ? ( n1597 ) : ( n1629 ) ;
assign n1631 =  ( n206 ) ? ( n1596 ) : ( n1630 ) ;
assign n1632 =  ( n205 ) ? ( n1595 ) : ( n1631 ) ;
assign n1633 =  ( n202 ) ? ( n1594 ) : ( n1632 ) ;
assign n1634 =  ( n199 ) ? ( n1593 ) : ( n1633 ) ;
assign n1635 =  ( n197 ) ? ( n1592 ) : ( n1634 ) ;
assign n1636 =  ( n195 ) ? ( n1591 ) : ( n1635 ) ;
assign n1637 =  ( n193 ) ? ( n1590 ) : ( n1636 ) ;
assign n1638 =  ( n191 ) ? ( n1589 ) : ( n1637 ) ;
assign n1639 =  ( n189 ) ? ( n1588 ) : ( n1638 ) ;
assign n1640 =  ( n187 ) ? ( n1587 ) : ( n1639 ) ;
assign n1641 =  ( n296 ) == ( 5'd30 )  ;
assign n1642 =  ( n1641 ) ? ( n300 ) : ( x30 ) ;
assign n1643 =  ( n1641 ) ? ( n302 ) : ( x30 ) ;
assign n1644 =  ( n1641 ) ? ( n304 ) : ( x30 ) ;
assign n1645 =  ( n1641 ) ? ( n306 ) : ( x30 ) ;
assign n1646 =  ( n1641 ) ? ( n308 ) : ( x30 ) ;
assign n1647 =  ( n1641 ) ? ( n310 ) : ( x30 ) ;
assign n1648 =  ( n1641 ) ? ( n312 ) : ( x30 ) ;
assign n1649 =  ( n1641 ) ? ( n314 ) : ( x30 ) ;
assign n1650 =  ( n1641 ) ? ( n316 ) : ( x30 ) ;
assign n1651 =  ( n1641 ) ? ( n318 ) : ( x30 ) ;
assign n1652 =  ( n1641 ) ? ( n321 ) : ( x30 ) ;
assign n1653 =  ( n1641 ) ? ( n323 ) : ( x30 ) ;
assign n1654 =  ( n1641 ) ? ( n325 ) : ( x30 ) ;
assign n1655 =  ( n1641 ) ? ( n328 ) : ( x30 ) ;
assign n1656 =  ( n1641 ) ? ( n439 ) : ( x30 ) ;
assign n1657 =  ( n1641 ) ? ( n333 ) : ( x30 ) ;
assign n1658 =  ( n1641 ) ? ( n553 ) : ( x30 ) ;
assign n1659 =  ( n1641 ) ? ( n339 ) : ( x30 ) ;
assign n1660 =  ( n1641 ) ? ( n341 ) : ( x30 ) ;
assign n1661 =  ( n1641 ) ? ( n162 ) : ( x30 ) ;
assign n1662 =  ( n1641 ) ? ( n347 ) : ( x30 ) ;
assign n1663 =  ( n1641 ) ? ( n346 ) : ( x30 ) ;
assign n1664 =  ( n1641 ) ? ( n370 ) : ( x30 ) ;
assign n1665 =  ( n1641 ) ? ( n378 ) : ( x30 ) ;
assign n1666 =  ( n1641 ) ? ( n387 ) : ( x30 ) ;
assign n1667 =  ( n1641 ) ? ( n393 ) : ( x30 ) ;
assign n1668 =  ( n1641 ) ? ( n395 ) : ( x30 ) ;
assign n1669 =  ( n230 ) ? ( n1668 ) : ( x30 ) ;
assign n1670 =  ( n229 ) ? ( n1667 ) : ( n1669 ) ;
assign n1671 =  ( n228 ) ? ( n1666 ) : ( n1670 ) ;
assign n1672 =  ( n227 ) ? ( n1665 ) : ( n1671 ) ;
assign n1673 =  ( n226 ) ? ( n1664 ) : ( n1672 ) ;
assign n1674 =  ( n220 ) ? ( n1663 ) : ( n1673 ) ;
assign n1675 =  ( n219 ) ? ( n1662 ) : ( n1674 ) ;
assign n1676 =  ( n343 ) ? ( n1661 ) : ( n1675 ) ;
assign n1677 =  ( n218 ) ? ( n1660 ) : ( n1676 ) ;
assign n1678 =  ( n217 ) ? ( n1659 ) : ( n1677 ) ;
assign n1679 =  ( n216 ) ? ( n1658 ) : ( n1678 ) ;
assign n1680 =  ( n215 ) ? ( n1657 ) : ( n1679 ) ;
assign n1681 =  ( n214 ) ? ( n1656 ) : ( n1680 ) ;
assign n1682 =  ( n213 ) ? ( n1655 ) : ( n1681 ) ;
assign n1683 =  ( n212 ) ? ( n1654 ) : ( n1682 ) ;
assign n1684 =  ( n210 ) ? ( n1653 ) : ( n1683 ) ;
assign n1685 =  ( n209 ) ? ( n1652 ) : ( n1684 ) ;
assign n1686 =  ( n206 ) ? ( n1651 ) : ( n1685 ) ;
assign n1687 =  ( n205 ) ? ( n1650 ) : ( n1686 ) ;
assign n1688 =  ( n202 ) ? ( n1649 ) : ( n1687 ) ;
assign n1689 =  ( n199 ) ? ( n1648 ) : ( n1688 ) ;
assign n1690 =  ( n197 ) ? ( n1647 ) : ( n1689 ) ;
assign n1691 =  ( n195 ) ? ( n1646 ) : ( n1690 ) ;
assign n1692 =  ( n193 ) ? ( n1645 ) : ( n1691 ) ;
assign n1693 =  ( n191 ) ? ( n1644 ) : ( n1692 ) ;
assign n1694 =  ( n189 ) ? ( n1643 ) : ( n1693 ) ;
assign n1695 =  ( n187 ) ? ( n1642 ) : ( n1694 ) ;
assign n1696 =  ( n296 ) == ( 5'd31 )  ;
assign n1697 =  ( n1696 ) ? ( n300 ) : ( x31 ) ;
assign n1698 =  ( n1696 ) ? ( n302 ) : ( x31 ) ;
assign n1699 =  ( n1696 ) ? ( n304 ) : ( x31 ) ;
assign n1700 =  ( n1696 ) ? ( n306 ) : ( x31 ) ;
assign n1701 =  ( n1696 ) ? ( n308 ) : ( x31 ) ;
assign n1702 =  ( n1696 ) ? ( n310 ) : ( x31 ) ;
assign n1703 =  ( n1696 ) ? ( n312 ) : ( x31 ) ;
assign n1704 =  ( n1696 ) ? ( n314 ) : ( x31 ) ;
assign n1705 =  ( n1696 ) ? ( n316 ) : ( x31 ) ;
assign n1706 =  ( n1696 ) ? ( n318 ) : ( x31 ) ;
assign n1707 =  ( n1696 ) ? ( n321 ) : ( x31 ) ;
assign n1708 =  ( n1696 ) ? ( n323 ) : ( x31 ) ;
assign n1709 =  ( n1696 ) ? ( n325 ) : ( x31 ) ;
assign n1710 =  ( n1696 ) ? ( n328 ) : ( x31 ) ;
assign n1711 =  ( n1696 ) ? ( n439 ) : ( x31 ) ;
assign n1712 =  ( n1696 ) ? ( n333 ) : ( x31 ) ;
assign n1713 =  ( n1696 ) ? ( n553 ) : ( x31 ) ;
assign n1714 =  ( n1696 ) ? ( n339 ) : ( x31 ) ;
assign n1715 =  ( n1696 ) ? ( n341 ) : ( x31 ) ;
assign n1716 =  ( n1696 ) ? ( n162 ) : ( x31 ) ;
assign n1717 =  ( n1696 ) ? ( n347 ) : ( x31 ) ;
assign n1718 =  ( n1696 ) ? ( n346 ) : ( x31 ) ;
assign n1719 =  ( n1696 ) ? ( n370 ) : ( x31 ) ;
assign n1720 =  ( n1696 ) ? ( n378 ) : ( x31 ) ;
assign n1721 =  ( n1696 ) ? ( n387 ) : ( x31 ) ;
assign n1722 =  ( n1696 ) ? ( n393 ) : ( x31 ) ;
assign n1723 =  ( n1696 ) ? ( n395 ) : ( x31 ) ;
assign n1724 =  ( n230 ) ? ( n1723 ) : ( x31 ) ;
assign n1725 =  ( n229 ) ? ( n1722 ) : ( n1724 ) ;
assign n1726 =  ( n228 ) ? ( n1721 ) : ( n1725 ) ;
assign n1727 =  ( n227 ) ? ( n1720 ) : ( n1726 ) ;
assign n1728 =  ( n226 ) ? ( n1719 ) : ( n1727 ) ;
assign n1729 =  ( n220 ) ? ( n1718 ) : ( n1728 ) ;
assign n1730 =  ( n219 ) ? ( n1717 ) : ( n1729 ) ;
assign n1731 =  ( n343 ) ? ( n1716 ) : ( n1730 ) ;
assign n1732 =  ( n218 ) ? ( n1715 ) : ( n1731 ) ;
assign n1733 =  ( n217 ) ? ( n1714 ) : ( n1732 ) ;
assign n1734 =  ( n216 ) ? ( n1713 ) : ( n1733 ) ;
assign n1735 =  ( n215 ) ? ( n1712 ) : ( n1734 ) ;
assign n1736 =  ( n214 ) ? ( n1711 ) : ( n1735 ) ;
assign n1737 =  ( n213 ) ? ( n1710 ) : ( n1736 ) ;
assign n1738 =  ( n212 ) ? ( n1709 ) : ( n1737 ) ;
assign n1739 =  ( n210 ) ? ( n1708 ) : ( n1738 ) ;
assign n1740 =  ( n209 ) ? ( n1707 ) : ( n1739 ) ;
assign n1741 =  ( n206 ) ? ( n1706 ) : ( n1740 ) ;
assign n1742 =  ( n205 ) ? ( n1705 ) : ( n1741 ) ;
assign n1743 =  ( n202 ) ? ( n1704 ) : ( n1742 ) ;
assign n1744 =  ( n199 ) ? ( n1703 ) : ( n1743 ) ;
assign n1745 =  ( n197 ) ? ( n1702 ) : ( n1744 ) ;
assign n1746 =  ( n195 ) ? ( n1701 ) : ( n1745 ) ;
assign n1747 =  ( n193 ) ? ( n1700 ) : ( n1746 ) ;
assign n1748 =  ( n191 ) ? ( n1699 ) : ( n1747 ) ;
assign n1749 =  ( n189 ) ? ( n1698 ) : ( n1748 ) ;
assign n1750 =  ( n187 ) ? ( n1697 ) : ( n1749 ) ;
assign n1751 =  ( n296 ) == ( 5'd4 )  ;
assign n1752 =  ( n1751 ) ? ( n300 ) : ( x4 ) ;
assign n1753 =  ( n1751 ) ? ( n302 ) : ( x4 ) ;
assign n1754 =  ( n1751 ) ? ( n304 ) : ( x4 ) ;
assign n1755 =  ( n1751 ) ? ( n306 ) : ( x4 ) ;
assign n1756 =  ( n1751 ) ? ( n308 ) : ( x4 ) ;
assign n1757 =  ( n1751 ) ? ( n310 ) : ( x4 ) ;
assign n1758 =  ( n1751 ) ? ( n312 ) : ( x4 ) ;
assign n1759 =  ( n1751 ) ? ( n314 ) : ( x4 ) ;
assign n1760 =  ( n1751 ) ? ( n316 ) : ( x4 ) ;
assign n1761 =  ( n1751 ) ? ( n318 ) : ( x4 ) ;
assign n1762 =  ( n1751 ) ? ( n321 ) : ( x4 ) ;
assign n1763 =  ( n1751 ) ? ( n323 ) : ( x4 ) ;
assign n1764 =  ( n1751 ) ? ( n325 ) : ( x4 ) ;
assign n1765 =  ( n1751 ) ? ( n328 ) : ( x4 ) ;
assign n1766 =  ( n1751 ) ? ( n439 ) : ( x4 ) ;
assign n1767 =  ( n1751 ) ? ( n333 ) : ( x4 ) ;
assign n1768 =  ( n1751 ) ? ( n553 ) : ( x4 ) ;
assign n1769 =  ( n1751 ) ? ( n339 ) : ( x4 ) ;
assign n1770 =  ( n1751 ) ? ( n341 ) : ( x4 ) ;
assign n1771 =  ( n1751 ) ? ( n162 ) : ( x4 ) ;
assign n1772 =  ( n1751 ) ? ( n347 ) : ( x4 ) ;
assign n1773 =  ( n1751 ) ? ( n346 ) : ( x4 ) ;
assign n1774 =  ( n1751 ) ? ( n370 ) : ( x4 ) ;
assign n1775 =  ( n1751 ) ? ( n378 ) : ( x4 ) ;
assign n1776 =  ( n1751 ) ? ( n387 ) : ( x4 ) ;
assign n1777 =  ( n1751 ) ? ( n393 ) : ( x4 ) ;
assign n1778 =  ( n1751 ) ? ( n395 ) : ( x4 ) ;
assign n1779 =  ( n230 ) ? ( n1778 ) : ( x4 ) ;
assign n1780 =  ( n229 ) ? ( n1777 ) : ( n1779 ) ;
assign n1781 =  ( n228 ) ? ( n1776 ) : ( n1780 ) ;
assign n1782 =  ( n227 ) ? ( n1775 ) : ( n1781 ) ;
assign n1783 =  ( n226 ) ? ( n1774 ) : ( n1782 ) ;
assign n1784 =  ( n220 ) ? ( n1773 ) : ( n1783 ) ;
assign n1785 =  ( n219 ) ? ( n1772 ) : ( n1784 ) ;
assign n1786 =  ( n343 ) ? ( n1771 ) : ( n1785 ) ;
assign n1787 =  ( n218 ) ? ( n1770 ) : ( n1786 ) ;
assign n1788 =  ( n217 ) ? ( n1769 ) : ( n1787 ) ;
assign n1789 =  ( n216 ) ? ( n1768 ) : ( n1788 ) ;
assign n1790 =  ( n215 ) ? ( n1767 ) : ( n1789 ) ;
assign n1791 =  ( n214 ) ? ( n1766 ) : ( n1790 ) ;
assign n1792 =  ( n213 ) ? ( n1765 ) : ( n1791 ) ;
assign n1793 =  ( n212 ) ? ( n1764 ) : ( n1792 ) ;
assign n1794 =  ( n210 ) ? ( n1763 ) : ( n1793 ) ;
assign n1795 =  ( n209 ) ? ( n1762 ) : ( n1794 ) ;
assign n1796 =  ( n206 ) ? ( n1761 ) : ( n1795 ) ;
assign n1797 =  ( n205 ) ? ( n1760 ) : ( n1796 ) ;
assign n1798 =  ( n202 ) ? ( n1759 ) : ( n1797 ) ;
assign n1799 =  ( n199 ) ? ( n1758 ) : ( n1798 ) ;
assign n1800 =  ( n197 ) ? ( n1757 ) : ( n1799 ) ;
assign n1801 =  ( n195 ) ? ( n1756 ) : ( n1800 ) ;
assign n1802 =  ( n193 ) ? ( n1755 ) : ( n1801 ) ;
assign n1803 =  ( n191 ) ? ( n1754 ) : ( n1802 ) ;
assign n1804 =  ( n189 ) ? ( n1753 ) : ( n1803 ) ;
assign n1805 =  ( n187 ) ? ( n1752 ) : ( n1804 ) ;
assign n1806 =  ( n296 ) == ( 5'd5 )  ;
assign n1807 =  ( n1806 ) ? ( n300 ) : ( x5 ) ;
assign n1808 =  ( n1806 ) ? ( n302 ) : ( x5 ) ;
assign n1809 =  ( n1806 ) ? ( n304 ) : ( x5 ) ;
assign n1810 =  ( n1806 ) ? ( n306 ) : ( x5 ) ;
assign n1811 =  ( n1806 ) ? ( n308 ) : ( x5 ) ;
assign n1812 =  ( n1806 ) ? ( n310 ) : ( x5 ) ;
assign n1813 =  ( n1806 ) ? ( n312 ) : ( x5 ) ;
assign n1814 =  ( n1806 ) ? ( n314 ) : ( x5 ) ;
assign n1815 =  ( n1806 ) ? ( n316 ) : ( x5 ) ;
assign n1816 =  ( n1806 ) ? ( n318 ) : ( x5 ) ;
assign n1817 =  ( n1806 ) ? ( n321 ) : ( x5 ) ;
assign n1818 =  ( n1806 ) ? ( n323 ) : ( x5 ) ;
assign n1819 =  ( n1806 ) ? ( n325 ) : ( x5 ) ;
assign n1820 =  ( n1806 ) ? ( n328 ) : ( x5 ) ;
assign n1821 =  ( n1806 ) ? ( n439 ) : ( x5 ) ;
assign n1822 =  ( n1806 ) ? ( n333 ) : ( x5 ) ;
assign n1823 =  ( n1806 ) ? ( n336 ) : ( x5 ) ;
assign n1824 =  ( n1806 ) ? ( n612 ) : ( x5 ) ;
assign n1825 =  ( n1806 ) ? ( n341 ) : ( x5 ) ;
assign n1826 =  ( n1806 ) ? ( n162 ) : ( x5 ) ;
assign n1827 =  ( n1806 ) ? ( n347 ) : ( x5 ) ;
assign n1828 =  ( n1806 ) ? ( n346 ) : ( x5 ) ;
assign n1829 =  ( n1806 ) ? ( n370 ) : ( x5 ) ;
assign n1830 =  ( n1806 ) ? ( n378 ) : ( x5 ) ;
assign n1831 =  ( n1806 ) ? ( n387 ) : ( x5 ) ;
assign n1832 =  ( n1806 ) ? ( n393 ) : ( x5 ) ;
assign n1833 =  ( n1806 ) ? ( n395 ) : ( x5 ) ;
assign n1834 =  ( n230 ) ? ( n1833 ) : ( x5 ) ;
assign n1835 =  ( n229 ) ? ( n1832 ) : ( n1834 ) ;
assign n1836 =  ( n228 ) ? ( n1831 ) : ( n1835 ) ;
assign n1837 =  ( n227 ) ? ( n1830 ) : ( n1836 ) ;
assign n1838 =  ( n226 ) ? ( n1829 ) : ( n1837 ) ;
assign n1839 =  ( n220 ) ? ( n1828 ) : ( n1838 ) ;
assign n1840 =  ( n219 ) ? ( n1827 ) : ( n1839 ) ;
assign n1841 =  ( n343 ) ? ( n1826 ) : ( n1840 ) ;
assign n1842 =  ( n218 ) ? ( n1825 ) : ( n1841 ) ;
assign n1843 =  ( n217 ) ? ( n1824 ) : ( n1842 ) ;
assign n1844 =  ( n216 ) ? ( n1823 ) : ( n1843 ) ;
assign n1845 =  ( n215 ) ? ( n1822 ) : ( n1844 ) ;
assign n1846 =  ( n214 ) ? ( n1821 ) : ( n1845 ) ;
assign n1847 =  ( n213 ) ? ( n1820 ) : ( n1846 ) ;
assign n1848 =  ( n212 ) ? ( n1819 ) : ( n1847 ) ;
assign n1849 =  ( n210 ) ? ( n1818 ) : ( n1848 ) ;
assign n1850 =  ( n209 ) ? ( n1817 ) : ( n1849 ) ;
assign n1851 =  ( n206 ) ? ( n1816 ) : ( n1850 ) ;
assign n1852 =  ( n205 ) ? ( n1815 ) : ( n1851 ) ;
assign n1853 =  ( n202 ) ? ( n1814 ) : ( n1852 ) ;
assign n1854 =  ( n199 ) ? ( n1813 ) : ( n1853 ) ;
assign n1855 =  ( n197 ) ? ( n1812 ) : ( n1854 ) ;
assign n1856 =  ( n195 ) ? ( n1811 ) : ( n1855 ) ;
assign n1857 =  ( n193 ) ? ( n1810 ) : ( n1856 ) ;
assign n1858 =  ( n191 ) ? ( n1809 ) : ( n1857 ) ;
assign n1859 =  ( n189 ) ? ( n1808 ) : ( n1858 ) ;
assign n1860 =  ( n187 ) ? ( n1807 ) : ( n1859 ) ;
assign n1861 =  ( n296 ) == ( 5'd6 )  ;
assign n1862 =  ( n1861 ) ? ( n300 ) : ( x6 ) ;
assign n1863 =  ( n1861 ) ? ( n302 ) : ( x6 ) ;
assign n1864 =  ( n1861 ) ? ( n304 ) : ( x6 ) ;
assign n1865 =  ( n1861 ) ? ( n306 ) : ( x6 ) ;
assign n1866 =  ( n1861 ) ? ( n308 ) : ( x6 ) ;
assign n1867 =  ( n1861 ) ? ( n310 ) : ( x6 ) ;
assign n1868 =  ( n1861 ) ? ( n312 ) : ( x6 ) ;
assign n1869 =  ( n1861 ) ? ( n314 ) : ( x6 ) ;
assign n1870 =  ( n1861 ) ? ( n316 ) : ( x6 ) ;
assign n1871 =  ( n1861 ) ? ( n318 ) : ( x6 ) ;
assign n1872 =  ( n1861 ) ? ( n321 ) : ( x6 ) ;
assign n1873 =  ( n1861 ) ? ( n323 ) : ( x6 ) ;
assign n1874 =  ( n1861 ) ? ( n325 ) : ( x6 ) ;
assign n1875 =  ( n1861 ) ? ( n328 ) : ( x6 ) ;
assign n1876 =  ( n1861 ) ? ( n439 ) : ( x6 ) ;
assign n1877 =  ( n1861 ) ? ( n333 ) : ( x6 ) ;
assign n1878 =  ( n1861 ) ? ( n553 ) : ( x6 ) ;
assign n1879 =  ( n1861 ) ? ( n339 ) : ( x6 ) ;
assign n1880 =  ( n70 ) + ( n330 )  ;
assign n1881 =  ( n1861 ) ? ( n1880 ) : ( x6 ) ;
assign n1882 =  ( n1861 ) ? ( n162 ) : ( x6 ) ;
assign n1883 =  ( n1861 ) ? ( n347 ) : ( x6 ) ;
assign n1884 =  ( n1861 ) ? ( n346 ) : ( x6 ) ;
assign n1885 =  ( n1861 ) ? ( n370 ) : ( x6 ) ;
assign n1886 =  ( n1861 ) ? ( n378 ) : ( x6 ) ;
assign n1887 =  ( n1861 ) ? ( n387 ) : ( x6 ) ;
assign n1888 =  ( n1861 ) ? ( n393 ) : ( x6 ) ;
assign n1889 =  ( n1861 ) ? ( n395 ) : ( x6 ) ;
assign n1890 =  ( n230 ) ? ( n1889 ) : ( x6 ) ;
assign n1891 =  ( n229 ) ? ( n1888 ) : ( n1890 ) ;
assign n1892 =  ( n228 ) ? ( n1887 ) : ( n1891 ) ;
assign n1893 =  ( n227 ) ? ( n1886 ) : ( n1892 ) ;
assign n1894 =  ( n226 ) ? ( n1885 ) : ( n1893 ) ;
assign n1895 =  ( n220 ) ? ( n1884 ) : ( n1894 ) ;
assign n1896 =  ( n219 ) ? ( n1883 ) : ( n1895 ) ;
assign n1897 =  ( n343 ) ? ( n1882 ) : ( n1896 ) ;
assign n1898 =  ( n218 ) ? ( n1881 ) : ( n1897 ) ;
assign n1899 =  ( n217 ) ? ( n1879 ) : ( n1898 ) ;
assign n1900 =  ( n216 ) ? ( n1878 ) : ( n1899 ) ;
assign n1901 =  ( n215 ) ? ( n1877 ) : ( n1900 ) ;
assign n1902 =  ( n214 ) ? ( n1876 ) : ( n1901 ) ;
assign n1903 =  ( n213 ) ? ( n1875 ) : ( n1902 ) ;
assign n1904 =  ( n212 ) ? ( n1874 ) : ( n1903 ) ;
assign n1905 =  ( n210 ) ? ( n1873 ) : ( n1904 ) ;
assign n1906 =  ( n209 ) ? ( n1872 ) : ( n1905 ) ;
assign n1907 =  ( n206 ) ? ( n1871 ) : ( n1906 ) ;
assign n1908 =  ( n205 ) ? ( n1870 ) : ( n1907 ) ;
assign n1909 =  ( n202 ) ? ( n1869 ) : ( n1908 ) ;
assign n1910 =  ( n199 ) ? ( n1868 ) : ( n1909 ) ;
assign n1911 =  ( n197 ) ? ( n1867 ) : ( n1910 ) ;
assign n1912 =  ( n195 ) ? ( n1866 ) : ( n1911 ) ;
assign n1913 =  ( n193 ) ? ( n1865 ) : ( n1912 ) ;
assign n1914 =  ( n191 ) ? ( n1864 ) : ( n1913 ) ;
assign n1915 =  ( n189 ) ? ( n1863 ) : ( n1914 ) ;
assign n1916 =  ( n187 ) ? ( n1862 ) : ( n1915 ) ;
assign n1917 =  ( n296 ) == ( 5'd7 )  ;
assign n1918 =  ( n1917 ) ? ( n300 ) : ( x7 ) ;
assign n1919 =  ( n1917 ) ? ( n302 ) : ( x7 ) ;
assign n1920 =  ( n1917 ) ? ( n304 ) : ( x7 ) ;
assign n1921 =  ( n1917 ) ? ( n306 ) : ( x7 ) ;
assign n1922 =  ( n1917 ) ? ( n308 ) : ( x7 ) ;
assign n1923 =  ( n1917 ) ? ( n310 ) : ( x7 ) ;
assign n1924 =  ( n1917 ) ? ( n312 ) : ( x7 ) ;
assign n1925 =  ( n1917 ) ? ( n314 ) : ( x7 ) ;
assign n1926 =  ( n1917 ) ? ( n316 ) : ( x7 ) ;
assign n1927 =  ( n1917 ) ? ( n318 ) : ( x7 ) ;
assign n1928 =  ( n1917 ) ? ( n321 ) : ( x7 ) ;
assign n1929 =  ( n1917 ) ? ( n323 ) : ( x7 ) ;
assign n1930 =  ( n1917 ) ? ( n325 ) : ( x7 ) ;
assign n1931 =  ( n1917 ) ? ( n328 ) : ( x7 ) ;
assign n1932 =  ( n1917 ) ? ( n439 ) : ( x7 ) ;
assign n1933 =  ( n1917 ) ? ( n333 ) : ( x7 ) ;
assign n1934 =  ( n1917 ) ? ( n553 ) : ( x7 ) ;
assign n1935 =  ( n1917 ) ? ( n339 ) : ( x7 ) ;
assign n1936 =  ( n1917 ) ? ( n341 ) : ( x7 ) ;
assign n1937 =  ( n1917 ) ? ( n162 ) : ( x7 ) ;
assign n1938 =  ( n1917 ) ? ( n347 ) : ( x7 ) ;
assign n1939 =  ( n1917 ) ? ( n346 ) : ( x7 ) ;
assign n1940 =  ( n1917 ) ? ( n370 ) : ( x7 ) ;
assign n1941 =  ( n1917 ) ? ( n378 ) : ( x7 ) ;
assign n1942 =  ( n1917 ) ? ( n387 ) : ( x7 ) ;
assign n1943 =  ( n1917 ) ? ( n393 ) : ( x7 ) ;
assign n1944 =  ( n1917 ) ? ( n395 ) : ( x7 ) ;
assign n1945 =  ( n230 ) ? ( n1944 ) : ( x7 ) ;
assign n1946 =  ( n229 ) ? ( n1943 ) : ( n1945 ) ;
assign n1947 =  ( n228 ) ? ( n1942 ) : ( n1946 ) ;
assign n1948 =  ( n227 ) ? ( n1941 ) : ( n1947 ) ;
assign n1949 =  ( n226 ) ? ( n1940 ) : ( n1948 ) ;
assign n1950 =  ( n220 ) ? ( n1939 ) : ( n1949 ) ;
assign n1951 =  ( n219 ) ? ( n1938 ) : ( n1950 ) ;
assign n1952 =  ( n343 ) ? ( n1937 ) : ( n1951 ) ;
assign n1953 =  ( n218 ) ? ( n1936 ) : ( n1952 ) ;
assign n1954 =  ( n217 ) ? ( n1935 ) : ( n1953 ) ;
assign n1955 =  ( n216 ) ? ( n1934 ) : ( n1954 ) ;
assign n1956 =  ( n215 ) ? ( n1933 ) : ( n1955 ) ;
assign n1957 =  ( n214 ) ? ( n1932 ) : ( n1956 ) ;
assign n1958 =  ( n213 ) ? ( n1931 ) : ( n1957 ) ;
assign n1959 =  ( n212 ) ? ( n1930 ) : ( n1958 ) ;
assign n1960 =  ( n210 ) ? ( n1929 ) : ( n1959 ) ;
assign n1961 =  ( n209 ) ? ( n1928 ) : ( n1960 ) ;
assign n1962 =  ( n206 ) ? ( n1927 ) : ( n1961 ) ;
assign n1963 =  ( n205 ) ? ( n1926 ) : ( n1962 ) ;
assign n1964 =  ( n202 ) ? ( n1925 ) : ( n1963 ) ;
assign n1965 =  ( n199 ) ? ( n1924 ) : ( n1964 ) ;
assign n1966 =  ( n197 ) ? ( n1923 ) : ( n1965 ) ;
assign n1967 =  ( n195 ) ? ( n1922 ) : ( n1966 ) ;
assign n1968 =  ( n193 ) ? ( n1921 ) : ( n1967 ) ;
assign n1969 =  ( n191 ) ? ( n1920 ) : ( n1968 ) ;
assign n1970 =  ( n189 ) ? ( n1919 ) : ( n1969 ) ;
assign n1971 =  ( n187 ) ? ( n1918 ) : ( n1970 ) ;
assign n1972 =  ( n296 ) == ( 5'd8 )  ;
assign n1973 =  ( n1972 ) ? ( n300 ) : ( x8 ) ;
assign n1974 =  ( n1972 ) ? ( n302 ) : ( x8 ) ;
assign n1975 =  ( n1972 ) ? ( n304 ) : ( x8 ) ;
assign n1976 =  ( n1972 ) ? ( n306 ) : ( x8 ) ;
assign n1977 =  ( n1972 ) ? ( n308 ) : ( x8 ) ;
assign n1978 =  ( n1972 ) ? ( n310 ) : ( x8 ) ;
assign n1979 =  ( n1972 ) ? ( n312 ) : ( x8 ) ;
assign n1980 =  ( n1972 ) ? ( n314 ) : ( x8 ) ;
assign n1981 =  ( n1972 ) ? ( n316 ) : ( x8 ) ;
assign n1982 =  ( n1972 ) ? ( n318 ) : ( x8 ) ;
assign n1983 =  ( n1972 ) ? ( n321 ) : ( x8 ) ;
assign n1984 =  ( n1972 ) ? ( n323 ) : ( x8 ) ;
assign n1985 =  ( n1972 ) ? ( n325 ) : ( x8 ) ;
assign n1986 =  ( n1972 ) ? ( n328 ) : ( x8 ) ;
assign n1987 =  ( n1972 ) ? ( n439 ) : ( x8 ) ;
assign n1988 =  ( n1972 ) ? ( n333 ) : ( x8 ) ;
assign n1989 =  ( n1972 ) ? ( n553 ) : ( x8 ) ;
assign n1990 =  ( n1972 ) ? ( n612 ) : ( x8 ) ;
assign n1991 =  ( n1972 ) ? ( n341 ) : ( x8 ) ;
assign n1992 =  ( n1972 ) ? ( n162 ) : ( x8 ) ;
assign n1993 =  ( n1972 ) ? ( n347 ) : ( x8 ) ;
assign n1994 =  ( n1972 ) ? ( n346 ) : ( x8 ) ;
assign n1995 =  ( n1972 ) ? ( n370 ) : ( x8 ) ;
assign n1996 =  ( n1972 ) ? ( n378 ) : ( x8 ) ;
assign n1997 =  ( n1972 ) ? ( n387 ) : ( x8 ) ;
assign n1998 =  ( n1972 ) ? ( n393 ) : ( x8 ) ;
assign n1999 =  ( n1972 ) ? ( n395 ) : ( x8 ) ;
assign n2000 =  ( n230 ) ? ( n1999 ) : ( x8 ) ;
assign n2001 =  ( n229 ) ? ( n1998 ) : ( n2000 ) ;
assign n2002 =  ( n228 ) ? ( n1997 ) : ( n2001 ) ;
assign n2003 =  ( n227 ) ? ( n1996 ) : ( n2002 ) ;
assign n2004 =  ( n226 ) ? ( n1995 ) : ( n2003 ) ;
assign n2005 =  ( n220 ) ? ( n1994 ) : ( n2004 ) ;
assign n2006 =  ( n219 ) ? ( n1993 ) : ( n2005 ) ;
assign n2007 =  ( n343 ) ? ( n1992 ) : ( n2006 ) ;
assign n2008 =  ( n218 ) ? ( n1991 ) : ( n2007 ) ;
assign n2009 =  ( n217 ) ? ( n1990 ) : ( n2008 ) ;
assign n2010 =  ( n216 ) ? ( n1989 ) : ( n2009 ) ;
assign n2011 =  ( n215 ) ? ( n1988 ) : ( n2010 ) ;
assign n2012 =  ( n214 ) ? ( n1987 ) : ( n2011 ) ;
assign n2013 =  ( n213 ) ? ( n1986 ) : ( n2012 ) ;
assign n2014 =  ( n212 ) ? ( n1985 ) : ( n2013 ) ;
assign n2015 =  ( n210 ) ? ( n1984 ) : ( n2014 ) ;
assign n2016 =  ( n209 ) ? ( n1983 ) : ( n2015 ) ;
assign n2017 =  ( n206 ) ? ( n1982 ) : ( n2016 ) ;
assign n2018 =  ( n205 ) ? ( n1981 ) : ( n2017 ) ;
assign n2019 =  ( n202 ) ? ( n1980 ) : ( n2018 ) ;
assign n2020 =  ( n199 ) ? ( n1979 ) : ( n2019 ) ;
assign n2021 =  ( n197 ) ? ( n1978 ) : ( n2020 ) ;
assign n2022 =  ( n195 ) ? ( n1977 ) : ( n2021 ) ;
assign n2023 =  ( n193 ) ? ( n1976 ) : ( n2022 ) ;
assign n2024 =  ( n191 ) ? ( n1975 ) : ( n2023 ) ;
assign n2025 =  ( n189 ) ? ( n1974 ) : ( n2024 ) ;
assign n2026 =  ( n187 ) ? ( n1973 ) : ( n2025 ) ;
assign n2027 =  ( n296 ) == ( 5'd9 )  ;
assign n2028 =  ( n2027 ) ? ( n300 ) : ( x9 ) ;
assign n2029 =  ( n2027 ) ? ( n302 ) : ( x9 ) ;
assign n2030 =  ( n2027 ) ? ( n304 ) : ( x9 ) ;
assign n2031 =  ( n2027 ) ? ( n306 ) : ( x9 ) ;
assign n2032 =  ( n2027 ) ? ( n308 ) : ( x9 ) ;
assign n2033 =  ( n2027 ) ? ( n310 ) : ( x9 ) ;
assign n2034 =  ( n2027 ) ? ( n312 ) : ( x9 ) ;
assign n2035 =  ( n2027 ) ? ( n314 ) : ( x9 ) ;
assign n2036 =  ( n2027 ) ? ( n316 ) : ( x9 ) ;
assign n2037 =  ( n2027 ) ? ( n318 ) : ( x9 ) ;
assign n2038 =  ( n2027 ) ? ( n321 ) : ( x9 ) ;
assign n2039 =  ( n2027 ) ? ( n323 ) : ( x9 ) ;
assign n2040 =  ( n2027 ) ? ( n325 ) : ( x9 ) ;
assign n2041 =  ( n2027 ) ? ( n719 ) : ( x9 ) ;
assign n2042 =  ( n2027 ) ? ( n439 ) : ( x9 ) ;
assign n2043 =  ( n2027 ) ? ( n333 ) : ( x9 ) ;
assign n2044 =  ( n2027 ) ? ( n553 ) : ( x9 ) ;
assign n2045 =  ( n2027 ) ? ( n612 ) : ( x9 ) ;
assign n2046 =  ( n2027 ) ? ( n341 ) : ( x9 ) ;
assign n2047 =  ( n2027 ) ? ( n162 ) : ( x9 ) ;
assign n2048 =  ( n2027 ) ? ( n347 ) : ( x9 ) ;
assign n2049 =  ( n2027 ) ? ( n346 ) : ( x9 ) ;
assign n2050 =  ( n2027 ) ? ( n370 ) : ( x9 ) ;
assign n2051 =  ( n2027 ) ? ( n378 ) : ( x9 ) ;
assign n2052 =  ( n2027 ) ? ( n387 ) : ( x9 ) ;
assign n2053 =  ( n2027 ) ? ( n393 ) : ( x9 ) ;
assign n2054 =  ( n2027 ) ? ( n395 ) : ( x9 ) ;
assign n2055 =  ( n230 ) ? ( n2054 ) : ( x9 ) ;
assign n2056 =  ( n229 ) ? ( n2053 ) : ( n2055 ) ;
assign n2057 =  ( n228 ) ? ( n2052 ) : ( n2056 ) ;
assign n2058 =  ( n227 ) ? ( n2051 ) : ( n2057 ) ;
assign n2059 =  ( n226 ) ? ( n2050 ) : ( n2058 ) ;
assign n2060 =  ( n220 ) ? ( n2049 ) : ( n2059 ) ;
assign n2061 =  ( n219 ) ? ( n2048 ) : ( n2060 ) ;
assign n2062 =  ( n343 ) ? ( n2047 ) : ( n2061 ) ;
assign n2063 =  ( n218 ) ? ( n2046 ) : ( n2062 ) ;
assign n2064 =  ( n217 ) ? ( n2045 ) : ( n2063 ) ;
assign n2065 =  ( n216 ) ? ( n2044 ) : ( n2064 ) ;
assign n2066 =  ( n215 ) ? ( n2043 ) : ( n2065 ) ;
assign n2067 =  ( n214 ) ? ( n2042 ) : ( n2066 ) ;
assign n2068 =  ( n213 ) ? ( n2041 ) : ( n2067 ) ;
assign n2069 =  ( n212 ) ? ( n2040 ) : ( n2068 ) ;
assign n2070 =  ( n210 ) ? ( n2039 ) : ( n2069 ) ;
assign n2071 =  ( n209 ) ? ( n2038 ) : ( n2070 ) ;
assign n2072 =  ( n206 ) ? ( n2037 ) : ( n2071 ) ;
assign n2073 =  ( n205 ) ? ( n2036 ) : ( n2072 ) ;
assign n2074 =  ( n202 ) ? ( n2035 ) : ( n2073 ) ;
assign n2075 =  ( n199 ) ? ( n2034 ) : ( n2074 ) ;
assign n2076 =  ( n197 ) ? ( n2033 ) : ( n2075 ) ;
assign n2077 =  ( n195 ) ? ( n2032 ) : ( n2076 ) ;
assign n2078 =  ( n193 ) ? ( n2031 ) : ( n2077 ) ;
assign n2079 =  ( n191 ) ? ( n2030 ) : ( n2078 ) ;
assign n2080 =  ( n189 ) ? ( n2029 ) : ( n2079 ) ;
assign n2081 =  ( n187 ) ? ( n2028 ) : ( n2080 ) ;
assign n2082 = ~ ( n222 ) ;
assign n2083 = ~ ( n223 ) ;
assign n2084 =  ( n2082 ) & ( n2083 )  ;
assign n2085 = ~ ( n224 ) ;
assign n2086 =  ( n2084 ) & ( n2085 )  ;
assign n2087 =  ( n2084 ) & ( n224 )  ;
assign n2088 =  { ( n185 ) , ( n296 ) }  ;
assign n2089 =  { {20{n2088[11] }  }, n2088}  ;
assign n2090 =  ( n70 ) + ( n2089 )  ;
assign n2091 = n2090[31:2] ;
assign n2092 =  {2'd0 , n2091}  ;
assign n2093 =  ( n151 ) & ( 32'd255 )  ;
assign n2094 = n2090[1:0] ;
assign n2095 =  {30'd0 , n2094}  ;
assign n2096 =  ( ( 32'd8 ) * ( n2095 ))  ;
assign n2097 =  ( n2093 ) << ( n2096 )  ;
assign n2098 =  ( 32'd255 ) << ( n2096 )  ;
assign n2099 = ~ ( n2098 ) ;
//assign n2100 =  (  mem [ n2092 ] )  ;
assign mem_raddr2 = n2092;
assign n2100 = mem_rdata2;

assign n2101 =  ( n2099 ) & ( n2100 )  ;
assign n2102 =  ( n2097 ) | ( n2101 )  ;
assign n2103 =  ( n2082 ) & ( n223 )  ;
assign n2104 =  ( n151 ) & ( 32'd65535 )  ;
assign n2105 =  ( n2104 ) << ( n2096 )  ;
assign n2106 =  ( 32'd65535 ) << ( n2096 )  ;
assign n2107 = ~ ( n2106 ) ;
assign n2108 =  ( n2107 ) & ( n2100 )  ;
assign n2109 =  ( n2105 ) | ( n2108 )  ;
assign n2110 =  ( n151 ) & ( 32'd4294967295 )  ;
assign n2111 =  ( n2110 ) << ( n2096 )  ;
assign n2112 =  ( 32'd4294967295 ) << ( n2096 )  ;
assign n2113 = ~ ( n2112 ) ;
assign n2114 =  ( n2113 ) & ( n2100 )  ;
assign n2115 =  ( n2111 ) | ( n2114 )  ;
assign mem_addr0 = n222 ? (n2092) : (n2103 ? (n2092) : (n2087 ? (n2092) : (0)));
assign mem_data0 = n222 ? (n2115) : (n2103 ? (n2109) : (n2087 ? (n2102) : (32'dx)));

assign mem_waddr0 = mem_addr0;
assign mem_wdata0 = mem_data0;
assign mem_wen0   = (n222 ? (1'b1) : (n2103 ? (1'b1) : (n2087 ? (1'b1) : (1'b0)))) & step;

always @(posedge clk) begin
   if(rst) begin
       pc <= pc;
       x0 <= x0;
       x1 <= x1;
       x10 <= x10;
       x11 <= x11;
       x12 <= x12;
       x13 <= x13;
       x14 <= x14;
       x15 <= x15;
       x16 <= x16;
       x17 <= x17;
       x18 <= x18;
       x19 <= x19;
       x2 <= x2;
       x20 <= x20;
       x21 <= x21;
       x22 <= x22;
       x23 <= x23;
       x24 <= x24;
       x25 <= x25;
       x26 <= x26;
       x27 <= x27;
       x28 <= x28;
       x29 <= x29;
       x3 <= x3;
       x30 <= x30;
       x31 <= x31;
       x4 <= x4;
       x5 <= x5;
       x6 <= x6;
       x7 <= x7;
       x8 <= x8;
       x9 <= x9;
   end
   else if(step) begin
       pc <= n267;
       x0 <= n295;
       x1 <= n423;
       x10 <= n479;
       x11 <= n534;
       x12 <= n591;
       x13 <= n649;
       x14 <= n704;
       x15 <= n760;
       x16 <= n815;
       x17 <= n870;
       x18 <= n925;
       x19 <= n980;
       x2 <= n1035;
       x20 <= n1090;
       x21 <= n1145;
       x22 <= n1200;
       x23 <= n1255;
       x24 <= n1310;
       x25 <= n1365;
       x26 <= n1420;
       x27 <= n1475;
       x28 <= n1530;
       x29 <= n1585;
       x3 <= n1640;
       x30 <= n1695;
       x31 <= n1750;
       x4 <= n1805;
       x5 <= n1860;
       x6 <= n1916;
       x7 <= n1971;
       x8 <= n2026;
       x9 <= n2081;
       //mem [ mem_addr0 ] <= mem_data0;
   end
end
endmodule
