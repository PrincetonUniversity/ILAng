module SPEC_B(
arg_0_TREADY,
arg_1_TDATA,
arg_1_TVALID,
LB1D_buff,
LB1D_in,
LB1D_it_1,
LB1D_p_cnt,
LB1D_uIn,
LB2D_proc_w,
LB2D_proc_x,
LB2D_proc_y,
LB2D_shift_0,
LB2D_shift_1,
LB2D_shift_2,
LB2D_shift_3,
LB2D_shift_4,
LB2D_shift_5,
LB2D_shift_6,
LB2D_shift_7,
LB2D_shift_x,
LB2D_shift_y,
arg_0_TDATA,
arg_0_TVALID,
arg_1_TREADY,
gb_exit_it_1,
gb_exit_it_2,
gb_exit_it_3,
gb_exit_it_4,
gb_exit_it_5,
gb_exit_it_6,
gb_exit_it_7,
gb_exit_it_8,
gb_p_cnt,
gb_pp_it_1,
gb_pp_it_2,
gb_pp_it_3,
gb_pp_it_4,
gb_pp_it_5,
gb_pp_it_6,
gb_pp_it_7,
gb_pp_it_8,
gb_pp_it_9,
in_stream_buff_0,
in_stream_buff_1,
in_stream_empty,
in_stream_full,
slice_stream_buff_0,
slice_stream_buff_1,
slice_stream_empty,
slice_stream_full,
stencil_stream_buff_0,
stencil_stream_buff_1,
stencil_stream_empty,
stencil_stream_full,
clk,rst,
step
);
input            arg_0_TREADY;
input      [7:0] arg_1_TDATA;
input            arg_1_TVALID;
input clk;
input rst;
input step;
output      [7:0] LB1D_buff;
output      [7:0] LB1D_in;
output            LB1D_it_1;
output     [18:0] LB1D_p_cnt;
output      [7:0] LB1D_uIn;
output     [63:0] LB2D_proc_w;
output      [8:0] LB2D_proc_x;
output      [9:0] LB2D_proc_y;
output     [71:0] LB2D_shift_0;
output     [71:0] LB2D_shift_1;
output     [71:0] LB2D_shift_2;
output     [71:0] LB2D_shift_3;
output     [71:0] LB2D_shift_4;
output     [71:0] LB2D_shift_5;
output     [71:0] LB2D_shift_6;
output     [71:0] LB2D_shift_7;
output      [8:0] LB2D_shift_x;
output      [9:0] LB2D_shift_y;
output      [7:0] arg_0_TDATA;
output            arg_0_TVALID;
output            arg_1_TREADY;
output            gb_exit_it_1;
output            gb_exit_it_2;
output            gb_exit_it_3;
output            gb_exit_it_4;
output            gb_exit_it_5;
output            gb_exit_it_6;
output            gb_exit_it_7;
output            gb_exit_it_8;
output     [18:0] gb_p_cnt;
output            gb_pp_it_1;
output            gb_pp_it_2;
output            gb_pp_it_3;
output            gb_pp_it_4;
output            gb_pp_it_5;
output            gb_pp_it_6;
output            gb_pp_it_7;
output            gb_pp_it_8;
output            gb_pp_it_9;
output      [7:0] in_stream_buff_0;
output      [7:0] in_stream_buff_1;
output            in_stream_empty;
output            in_stream_full;
output     [71:0] slice_stream_buff_0;
output     [71:0] slice_stream_buff_1;
output            slice_stream_empty;
output            slice_stream_full;
output    [647:0] stencil_stream_buff_0;
output    [647:0] stencil_stream_buff_1;
output            stencil_stream_empty;
output            stencil_stream_full;
reg      [7:0] LB1D_buff;
reg      [7:0] LB1D_in;
reg            LB1D_it_1;
reg     [18:0] LB1D_p_cnt;
reg      [7:0] LB1D_uIn;
reg     [63:0] LB2D_proc_w;
reg      [8:0] LB2D_proc_x;
reg      [9:0] LB2D_proc_y;
reg     [71:0] LB2D_shift_0;
reg     [71:0] LB2D_shift_1;
reg     [71:0] LB2D_shift_2;
reg     [71:0] LB2D_shift_3;
reg     [71:0] LB2D_shift_4;
reg     [71:0] LB2D_shift_5;
reg     [71:0] LB2D_shift_6;
reg     [71:0] LB2D_shift_7;
reg      [8:0] LB2D_shift_x;
reg      [9:0] LB2D_shift_y;
reg      [7:0] arg_0_TDATA;
reg            arg_0_TVALID;
reg            arg_1_TREADY;
reg            gb_exit_it_1;
reg            gb_exit_it_2;
reg            gb_exit_it_3;
reg            gb_exit_it_4;
reg            gb_exit_it_5;
reg            gb_exit_it_6;
reg            gb_exit_it_7;
reg            gb_exit_it_8;
reg     [18:0] gb_p_cnt;
reg            gb_pp_it_1;
reg            gb_pp_it_2;
reg            gb_pp_it_3;
reg            gb_pp_it_4;
reg            gb_pp_it_5;
reg            gb_pp_it_6;
reg            gb_pp_it_7;
reg            gb_pp_it_8;
reg            gb_pp_it_9;
reg      [7:0] in_stream_buff_0;
reg      [7:0] in_stream_buff_1;
reg            in_stream_empty;
reg            in_stream_full;
reg     [71:0] slice_stream_buff_0;
reg     [71:0] slice_stream_buff_1;
reg            slice_stream_empty;
reg            slice_stream_full;
reg    [647:0] stencil_stream_buff_0;
reg    [647:0] stencil_stream_buff_1;
reg            stencil_stream_empty;
reg            stencil_stream_full;
wire            arg_0_TREADY;
wire      [7:0] arg_1_TDATA;
wire            arg_1_TVALID;
wire            n0;
wire            n1;
wire            n2;
wire            n3;
wire            n4;
wire            n5;
wire            n6;
wire            n7;
wire            n8;
wire            n9;
wire            n10;
wire            n11;
wire            n12;
wire            n13;
wire            n14;
wire            n15;
wire            n16;
wire            n17;
wire            n18;
wire            n19;
wire            n20;
wire            n21;
wire            n22;
wire            n23;
wire            n24;
wire            n25;
wire            n26;
wire            n27;
wire            n28;
wire            n29;
wire            n30;
wire            n31;
wire            n32;
wire            n33;
wire            n34;
wire            n35;
wire            n36;
wire            n37;
wire            n38;
wire      [7:0] n39;
wire      [7:0] n40;
wire      [7:0] n41;
wire      [7:0] n42;
wire      [7:0] n43;
wire      [7:0] n44;
wire      [7:0] n45;
wire      [7:0] n46;
wire      [7:0] n47;
wire      [7:0] n48;
wire      [7:0] n49;
wire      [7:0] n50;
wire      [7:0] n51;
wire      [7:0] n52;
wire            n53;
wire            n54;
wire            n55;
wire     [18:0] n56;
wire     [18:0] n57;
wire     [18:0] n58;
wire     [18:0] n59;
wire     [18:0] n60;
wire     [18:0] n61;
wire     [18:0] n62;
wire     [18:0] n63;
wire      [7:0] n64;
wire      [7:0] n65;
wire      [7:0] n66;
wire      [7:0] n67;
wire      [7:0] n68;
wire      [7:0] n69;
wire      [7:0] n70;
wire            n71;
wire            n72;
wire     [63:0] n73;
wire     [63:0] n74;
wire     [63:0] n75;
wire     [63:0] n76;
wire     [63:0] n77;
wire     [63:0] n78;
wire     [63:0] n79;
wire     [63:0] n80;
wire      [8:0] n81;
wire      [8:0] n82;
wire      [8:0] n83;
wire      [8:0] n84;
wire      [8:0] n85;
wire      [8:0] n86;
wire      [8:0] n87;
wire            n88;
wire      [9:0] n89;
wire      [9:0] n90;
wire      [9:0] n91;
wire      [9:0] n92;
wire      [9:0] n93;
wire      [9:0] n94;
wire      [9:0] n95;
wire      [9:0] n96;
wire     [71:0] n97;
wire     [71:0] n98;
wire     [71:0] n99;
wire     [71:0] n100;
wire     [71:0] n101;
wire     [71:0] n102;
wire     [71:0] n103;
wire     [71:0] n104;
wire     [71:0] n105;
wire     [71:0] n106;
wire     [71:0] n107;
wire     [71:0] n108;
wire     [71:0] n109;
wire     [71:0] n110;
wire     [71:0] n111;
wire     [71:0] n112;
wire     [71:0] n113;
wire     [71:0] n114;
wire     [71:0] n115;
wire     [71:0] n116;
wire     [71:0] n117;
wire     [71:0] n118;
wire     [71:0] n119;
wire     [71:0] n120;
wire     [71:0] n121;
wire     [71:0] n122;
wire     [71:0] n123;
wire     [71:0] n124;
wire     [71:0] n125;
wire     [71:0] n126;
wire     [71:0] n127;
wire     [71:0] n128;
wire     [71:0] n129;
wire     [71:0] n130;
wire     [71:0] n131;
wire            n132;
wire     [71:0] n133;
wire     [71:0] n134;
wire     [71:0] n135;
wire     [71:0] n136;
wire     [71:0] n137;
wire     [71:0] n138;
wire            n139;
wire            n140;
wire            n141;
wire            n142;
wire      [8:0] n143;
wire      [8:0] n144;
wire      [8:0] n145;
wire      [8:0] n146;
wire      [8:0] n147;
wire      [8:0] n148;
wire      [8:0] n149;
wire            n150;
wire            n151;
wire      [9:0] n152;
wire      [9:0] n153;
wire      [9:0] n154;
wire      [9:0] n155;
wire      [9:0] n156;
wire      [9:0] n157;
wire      [9:0] n158;
wire      [9:0] n159;
wire            n160;
wire    [647:0] n161;
wire      [7:0] n162;
wire      [7:0] n163;
wire      [7:0] n164;
wire      [7:0] n165;
wire      [7:0] n166;
wire      [7:0] n167;
wire      [7:0] n168;
wire            n169;
wire            n170;
wire            n171;
wire            n172;
wire            n173;
wire            n174;
wire            n175;
wire            n176;
wire            n177;
wire            n178;
wire            n179;
wire            n180;
wire            n181;
wire            n182;
wire            n183;
wire     [18:0] n184;
wire            n185;
wire            n186;
wire            n187;
wire            n188;
wire            n189;
wire            n190;
wire            n191;
wire            n192;
wire            n193;
wire            n194;
wire            n195;
wire            n196;
wire            n197;
wire            n198;
wire            n199;
wire            n200;
wire            n201;
wire            n202;
wire            n203;
wire            n204;
wire            n205;
wire            n206;
wire            n207;
wire            n208;
wire            n209;
wire            n210;
wire            n211;
wire            n212;
wire            n213;
wire            n214;
wire            n215;
wire            n216;
wire            n217;
wire            n218;
wire            n219;
wire            n220;
wire            n221;
wire            n222;
wire            n223;
wire            n224;
wire            n225;
wire            n226;
wire            n227;
wire     [18:0] n228;
wire     [18:0] n229;
wire     [18:0] n230;
wire     [18:0] n231;
wire     [18:0] n232;
wire     [18:0] n233;
wire            n234;
wire            n235;
wire            n236;
wire            n237;
wire            n238;
wire            n239;
wire            n240;
wire            n241;
wire            n242;
wire            n243;
wire            n244;
wire            n245;
wire            n246;
wire            n247;
wire            n248;
wire            n249;
wire            n250;
wire            n251;
wire            n252;
wire            n253;
wire            n254;
wire            n255;
wire            n256;
wire            n257;
wire            n258;
wire            n259;
wire            n260;
wire            n261;
wire            n262;
wire            n263;
wire            n264;
wire            n265;
wire            n266;
wire            n267;
wire            n268;
wire            n269;
wire            n270;
wire            n271;
wire            n272;
wire            n273;
wire            n274;
wire            n275;
wire            n276;
wire            n277;
wire            n278;
wire      [7:0] n279;
wire      [7:0] n280;
wire      [7:0] n281;
wire      [7:0] n282;
wire      [7:0] n283;
wire      [7:0] n284;
wire      [7:0] n285;
wire      [7:0] n286;
wire      [7:0] n287;
wire      [7:0] n288;
wire      [7:0] n289;
wire      [7:0] n290;
wire            n291;
wire            n292;
wire            n293;
wire            n294;
wire            n295;
wire            n296;
wire            n297;
wire            n298;
wire            n299;
wire            n300;
wire            n301;
wire            n302;
wire            n303;
wire            n304;
wire            n305;
wire            n306;
wire      [7:0] n307;
wire            n308;
wire      [8:0] n309;
wire      [7:0] n310;
wire            n311;
wire      [7:0] n312;
wire            n313;
wire      [7:0] n314;
wire            n315;
wire      [7:0] n316;
wire            n317;
wire      [7:0] n318;
wire            n319;
wire      [7:0] n320;
wire            n321;
wire      [7:0] n322;
wire      [7:0] n323;
wire      [7:0] n324;
wire      [7:0] n325;
wire      [7:0] n326;
wire      [7:0] n327;
wire      [7:0] n328;
wire      [7:0] n329;
wire      [7:0] n330;
wire      [7:0] n331;
wire      [7:0] n332;
wire      [7:0] n333;
wire      [7:0] n334;
wire      [7:0] n335;
wire      [7:0] n336;
wire      [7:0] n337;
wire      [7:0] n338;
wire      [7:0] n339;
wire      [7:0] n340;
wire      [7:0] n341;
wire      [7:0] n342;
wire      [7:0] n343;
wire      [7:0] n344;
wire      [7:0] n345;
wire      [7:0] n346;
wire      [7:0] n347;
wire      [7:0] n348;
wire      [7:0] n349;
wire      [7:0] n350;
wire      [7:0] n351;
wire      [7:0] n352;
wire      [7:0] n353;
wire      [7:0] n354;
wire      [7:0] n355;
wire      [7:0] n356;
wire      [7:0] n357;
wire      [7:0] n358;
wire      [7:0] n359;
wire      [7:0] n360;
wire      [7:0] n361;
wire      [7:0] n362;
wire      [7:0] n363;
wire      [7:0] n364;
wire      [7:0] n365;
wire      [7:0] n366;
wire      [7:0] n367;
wire      [7:0] n368;
wire      [7:0] n369;
wire      [7:0] n370;
wire      [7:0] n371;
wire      [7:0] n372;
wire      [7:0] n373;
wire      [7:0] n374;
wire      [7:0] n375;
wire      [7:0] n376;
wire      [7:0] n377;
wire      [7:0] n378;
wire      [7:0] n379;
wire     [15:0] n380;
wire     [23:0] n381;
wire     [31:0] n382;
wire     [39:0] n383;
wire     [47:0] n384;
wire     [55:0] n385;
wire     [63:0] n386;
wire     [71:0] n387;
wire     [71:0] n388;
wire     [71:0] n389;
wire     [71:0] n390;
wire     [71:0] n391;
wire     [71:0] n392;
wire     [71:0] n393;
wire     [71:0] n394;
wire     [71:0] n395;
wire     [71:0] n396;
wire     [71:0] n397;
wire     [71:0] n398;
wire     [71:0] n399;
wire            n400;
wire            n401;
wire            n402;
wire            n403;
wire            n404;
wire            n405;
wire            n406;
wire            n407;
wire            n408;
wire            n409;
wire            n410;
wire            n411;
wire            n412;
wire            n413;
wire            n414;
wire            n415;
wire            n416;
wire            n417;
wire      [7:0] n418;
wire      [7:0] n419;
wire      [7:0] n420;
wire      [7:0] n421;
wire      [7:0] n422;
wire      [7:0] n423;
wire      [7:0] n424;
wire      [7:0] n425;
wire      [7:0] n426;
wire     [15:0] n427;
wire     [23:0] n428;
wire     [31:0] n429;
wire     [39:0] n430;
wire     [47:0] n431;
wire     [55:0] n432;
wire     [63:0] n433;
wire     [71:0] n434;
wire      [7:0] n435;
wire      [7:0] n436;
wire      [7:0] n437;
wire      [7:0] n438;
wire      [7:0] n439;
wire      [7:0] n440;
wire      [7:0] n441;
wire      [7:0] n442;
wire      [7:0] n443;
wire     [15:0] n444;
wire     [23:0] n445;
wire     [31:0] n446;
wire     [39:0] n447;
wire     [47:0] n448;
wire     [55:0] n449;
wire     [63:0] n450;
wire     [71:0] n451;
wire      [7:0] n452;
wire      [7:0] n453;
wire      [7:0] n454;
wire      [7:0] n455;
wire      [7:0] n456;
wire      [7:0] n457;
wire      [7:0] n458;
wire      [7:0] n459;
wire      [7:0] n460;
wire     [15:0] n461;
wire     [23:0] n462;
wire     [31:0] n463;
wire     [39:0] n464;
wire     [47:0] n465;
wire     [55:0] n466;
wire     [63:0] n467;
wire     [71:0] n468;
wire      [7:0] n469;
wire      [7:0] n470;
wire      [7:0] n471;
wire      [7:0] n472;
wire      [7:0] n473;
wire      [7:0] n474;
wire      [7:0] n475;
wire      [7:0] n476;
wire      [7:0] n477;
wire     [15:0] n478;
wire     [23:0] n479;
wire     [31:0] n480;
wire     [39:0] n481;
wire     [47:0] n482;
wire     [55:0] n483;
wire     [63:0] n484;
wire     [71:0] n485;
wire      [7:0] n486;
wire      [7:0] n487;
wire      [7:0] n488;
wire      [7:0] n489;
wire      [7:0] n490;
wire      [7:0] n491;
wire      [7:0] n492;
wire      [7:0] n493;
wire      [7:0] n494;
wire     [15:0] n495;
wire     [23:0] n496;
wire     [31:0] n497;
wire     [39:0] n498;
wire     [47:0] n499;
wire     [55:0] n500;
wire     [63:0] n501;
wire     [71:0] n502;
wire      [7:0] n503;
wire      [7:0] n504;
wire      [7:0] n505;
wire      [7:0] n506;
wire      [7:0] n507;
wire      [7:0] n508;
wire      [7:0] n509;
wire      [7:0] n510;
wire      [7:0] n511;
wire     [15:0] n512;
wire     [23:0] n513;
wire     [31:0] n514;
wire     [39:0] n515;
wire     [47:0] n516;
wire     [55:0] n517;
wire     [63:0] n518;
wire     [71:0] n519;
wire      [7:0] n520;
wire      [7:0] n521;
wire      [7:0] n522;
wire      [7:0] n523;
wire      [7:0] n524;
wire      [7:0] n525;
wire      [7:0] n526;
wire      [7:0] n527;
wire      [7:0] n528;
wire     [15:0] n529;
wire     [23:0] n530;
wire     [31:0] n531;
wire     [39:0] n532;
wire     [47:0] n533;
wire     [55:0] n534;
wire     [63:0] n535;
wire     [71:0] n536;
wire      [7:0] n537;
wire      [7:0] n538;
wire      [7:0] n539;
wire      [7:0] n540;
wire      [7:0] n541;
wire      [7:0] n542;
wire      [7:0] n543;
wire      [7:0] n544;
wire      [7:0] n545;
wire     [15:0] n546;
wire     [23:0] n547;
wire     [31:0] n548;
wire     [39:0] n549;
wire     [47:0] n550;
wire     [55:0] n551;
wire     [63:0] n552;
wire     [71:0] n553;
wire      [7:0] n554;
wire      [7:0] n555;
wire      [7:0] n556;
wire      [7:0] n557;
wire      [7:0] n558;
wire      [7:0] n559;
wire      [7:0] n560;
wire      [7:0] n561;
wire      [7:0] n562;
wire     [15:0] n563;
wire     [23:0] n564;
wire     [31:0] n565;
wire     [39:0] n566;
wire     [47:0] n567;
wire     [55:0] n568;
wire     [63:0] n569;
wire     [71:0] n570;
wire    [143:0] n571;
wire    [215:0] n572;
wire    [287:0] n573;
wire    [359:0] n574;
wire    [431:0] n575;
wire    [503:0] n576;
wire    [575:0] n577;
wire    [647:0] n578;
wire    [647:0] n579;
wire    [647:0] n580;
wire    [647:0] n581;
wire    [647:0] n582;
wire    [647:0] n583;
wire    [647:0] n584;
wire    [647:0] n585;
wire    [647:0] n586;
wire    [647:0] n587;
wire    [647:0] n588;
wire    [647:0] n589;
wire            n590;
wire            n591;
wire            n592;
wire            n593;
wire            n594;
wire            n595;
wire            n596;
wire            n597;
wire            n598;
wire            n599;
wire            n600;
wire            n601;
wire            n602;
wire            n603;
wire            n604;
wire            n605;
wire            n606;
wire      [8:0] LB2D_proc_0_addr0;
wire      [7:0] LB2D_proc_0_data0;
wire            n607;
wire            n608;
wire            n609;
wire            n610;
wire            n611;
wire            n612;
wire            n613;
wire            n614;
wire            n615;
wire            n616;
wire            n617;
wire            n618;
wire            n619;
wire            n620;
wire            n621;
wire            n622;
wire      [8:0] LB2D_proc_1_addr0;
wire      [7:0] LB2D_proc_1_data0;
wire            n623;
wire            n624;
wire            n625;
wire      [8:0] LB2D_proc_2_addr0;
wire      [7:0] LB2D_proc_2_data0;
wire            n626;
wire            n627;
wire            n628;
wire      [8:0] LB2D_proc_3_addr0;
wire      [7:0] LB2D_proc_3_data0;
wire            n629;
wire            n630;
wire            n631;
wire      [8:0] LB2D_proc_4_addr0;
wire      [7:0] LB2D_proc_4_data0;
wire            n632;
wire            n633;
wire            n634;
wire      [8:0] LB2D_proc_5_addr0;
wire      [7:0] LB2D_proc_5_data0;
wire            n635;
wire            n636;
wire            n637;
wire      [8:0] LB2D_proc_6_addr0;
wire      [7:0] LB2D_proc_6_data0;
wire            n638;
wire            n639;
wire            n640;
wire      [8:0] LB2D_proc_7_addr0;
wire      [7:0] LB2D_proc_7_data0;
wire            n641;
wire            n642;
wire            n643;
reg      [7:0] LB2D_proc_0[511:0];
reg      [7:0] LB2D_proc_1[511:0];
reg      [7:0] LB2D_proc_2[511:0];
reg      [7:0] LB2D_proc_3[511:0];
reg      [7:0] LB2D_proc_4[511:0];
reg      [7:0] LB2D_proc_5[511:0];
reg      [7:0] LB2D_proc_6[511:0];
reg      [7:0] LB2D_proc_7[511:0];
wire clk;
wire rst;
wire step;
assign n0 =  ( arg_1_TREADY ) == ( 1'd1 )  ;
assign n1 =  ( arg_1_TVALID ) == ( 1'd1 )  ;
assign n2 =  ( n0 ) & ( n1 )  ;
assign n3 =  ( arg_0_TREADY ) == ( 1'd0 )  ;
assign n4 =  ( n2 ) & ( n3 )  ;
assign n5 =  ( arg_0_TVALID ) == ( 1'd0 )  ;
assign n6 =  ( gb_exit_it_1 ) == ( 1'd0 )  ;
assign n7 =  ( stencil_stream_empty ) == ( 1'd0 )  ;
assign n8 =  ( n6 ) & ( n7 )  ;
assign n9 =  ( gb_exit_it_1 ) == ( 1'd1 )  ;
assign n10 =  ( gb_exit_it_8 ) == ( 1'd0 )  ;
assign n11 =  ( n9 ) & ( n10 )  ;
assign n12 =  ( n8 ) | ( n11 )  ;
assign n13 =  ( n5 ) & ( n12 )  ;
assign n14 =  ( slice_stream_empty ) == ( 1'd0 )  ;
assign n15 =  ( LB2D_shift_x ) != ( 9'd488 )  ;
assign n16 =  ( n14 ) & ( n15 )  ;
assign n17 =  ( stencil_stream_full ) == ( 1'd0 )  ;
assign n18 =  ( LB2D_shift_x ) < ( 9'd8 )  ;
assign n19 =  ( LB2D_shift_x ) > ( 9'd0 )  ;
assign n20 =  ( n18 ) & ( n19 )  ;
assign n21 =  ( n17 ) | ( n20 )  ;
assign n22 =  ( n16 ) & ( n21 )  ;
assign n23 =  ( in_stream_empty ) == ( 1'd0 )  ;
assign n24 =  ( slice_stream_full ) == ( 1'd0 )  ;
assign n25 =  ( LB2D_proc_y ) < ( 10'd8 )  ;
assign n26 =  ( n24 ) | ( n25 )  ;
assign n27 =  ( n23 ) & ( n26 )  ;
assign n28 =  ( in_stream_full ) == ( 1'd0 )  ;
assign n29 =  ( n0 ) & ( n28 )  ;
assign n30 =  ( LB1D_it_1 ) == ( 1'd1 )  ;
assign n31 =  ( n29 ) & ( n30 )  ;
assign n32 =  ( LB1D_p_cnt ) == ( 19'd316224 )  ;
assign n33 =  ( n31 ) & ( n32 )  ;
assign n34 =  ( arg_1_TREADY ) == ( 1'd0 )  ;
assign n35 =  ( n34 ) & ( n28 )  ;
assign n36 =  ( LB1D_it_1 ) == ( 1'd0 )  ;
assign n37 =  ( n35 ) & ( n36 )  ;
assign n38 =  ( n35 ) & ( n30 )  ;
assign n39 =  ( n38 ) ? ( LB1D_uIn ) : ( LB1D_buff ) ;
assign n40 =  ( n37 ) ? ( LB1D_uIn ) : ( n39 ) ;
assign n41 =  ( n33 ) ? ( LB1D_uIn ) : ( n40 ) ;
assign n42 =  ( n27 ) ? ( LB1D_buff ) : ( n41 ) ;
assign n43 =  ( n22 ) ? ( LB1D_buff ) : ( n42 ) ;
assign n44 =  ( n13 ) ? ( LB1D_buff ) : ( n43 ) ;
assign n45 =  ( n4 ) ? ( LB1D_buff ) : ( n44 ) ;
assign n46 =  ( n38 ) ? ( LB1D_in ) : ( LB1D_in ) ;
assign n47 =  ( n37 ) ? ( LB1D_in ) : ( n46 ) ;
assign n48 =  ( n33 ) ? ( LB1D_in ) : ( n47 ) ;
assign n49 =  ( n27 ) ? ( LB1D_in ) : ( n48 ) ;
assign n50 =  ( n22 ) ? ( LB1D_in ) : ( n49 ) ;
assign n51 =  ( n13 ) ? ( LB1D_in ) : ( n50 ) ;
assign n52 =  ( n4 ) ? ( arg_1_TDATA ) : ( n51 ) ;
assign n53 =  ( n38 ) ? ( 1'd1 ) : ( LB1D_it_1 ) ;
assign n54 =  ( n37 ) ? ( 1'd1 ) : ( n53 ) ;
assign n55 =  ( n33 ) ? ( 1'd0 ) : ( n54 ) ;
assign n56 =  ( LB1D_p_cnt ) + ( 19'd1 )  ;
assign n57 =  ( n38 ) ? ( n56 ) : ( LB1D_p_cnt ) ;
assign n58 =  ( n37 ) ? ( n56 ) : ( n57 ) ;
assign n59 =  ( n33 ) ? ( 19'd0 ) : ( n58 ) ;
assign n60 =  ( n27 ) ? ( LB1D_p_cnt ) : ( n59 ) ;
assign n61 =  ( n22 ) ? ( LB1D_p_cnt ) : ( n60 ) ;
assign n62 =  ( n13 ) ? ( LB1D_p_cnt ) : ( n61 ) ;
assign n63 =  ( n4 ) ? ( LB1D_p_cnt ) : ( n62 ) ;
assign n64 =  ( n38 ) ? ( LB1D_in ) : ( LB1D_uIn ) ;
assign n65 =  ( n37 ) ? ( LB1D_in ) : ( n64 ) ;
assign n66 =  ( n33 ) ? ( LB1D_in ) : ( n65 ) ;
assign n67 =  ( n27 ) ? ( LB1D_uIn ) : ( n66 ) ;
assign n68 =  ( n22 ) ? ( LB1D_uIn ) : ( n67 ) ;
assign n69 =  ( n13 ) ? ( LB1D_uIn ) : ( n68 ) ;
assign n70 =  ( n4 ) ? ( LB1D_uIn ) : ( n69 ) ;
assign n71 =  ( LB2D_proc_x ) == ( 9'd488 )  ;
assign n72 =  ( LB2D_proc_w ) == ( 64'd7 )  ;
assign n73 =  ( LB2D_proc_w ) + ( 64'd1 )  ;
assign n74 =  ( n72 ) ? ( 64'd0 ) : ( n73 ) ;
assign n75 =  ( n71 ) ? ( n74 ) : ( LB2D_proc_w ) ;
assign n76 =  ( n38 ) ? ( LB2D_proc_w ) : ( LB2D_proc_w ) ;
assign n77 =  ( n27 ) ? ( n75 ) : ( n76 ) ;
assign n78 =  ( n22 ) ? ( LB2D_proc_w ) : ( n77 ) ;
assign n79 =  ( n13 ) ? ( LB2D_proc_w ) : ( n78 ) ;
assign n80 =  ( n4 ) ? ( LB2D_proc_w ) : ( n79 ) ;
assign n81 =  ( LB2D_proc_x ) + ( 9'd1 )  ;
assign n82 =  ( n71 ) ? ( 9'd1 ) : ( n81 ) ;
assign n83 =  ( n38 ) ? ( LB2D_proc_x ) : ( LB2D_proc_x ) ;
assign n84 =  ( n27 ) ? ( n82 ) : ( n83 ) ;
assign n85 =  ( n22 ) ? ( LB2D_proc_x ) : ( n84 ) ;
assign n86 =  ( n13 ) ? ( LB2D_proc_x ) : ( n85 ) ;
assign n87 =  ( n4 ) ? ( LB2D_proc_x ) : ( n86 ) ;
assign n88 =  ( LB2D_proc_y ) == ( 10'd648 )  ;
assign n89 =  ( LB2D_proc_y ) + ( 10'd1 )  ;
assign n90 =  ( n88 ) ? ( 10'd0 ) : ( n89 ) ;
assign n91 =  ( n71 ) ? ( n90 ) : ( LB2D_proc_y ) ;
assign n92 =  ( n38 ) ? ( LB2D_proc_y ) : ( LB2D_proc_y ) ;
assign n93 =  ( n27 ) ? ( n91 ) : ( n92 ) ;
assign n94 =  ( n22 ) ? ( LB2D_proc_y ) : ( n93 ) ;
assign n95 =  ( n13 ) ? ( LB2D_proc_y ) : ( n94 ) ;
assign n96 =  ( n4 ) ? ( LB2D_proc_y ) : ( n95 ) ;
assign n97 =  ( n38 ) ? ( LB2D_shift_0 ) : ( LB2D_shift_0 ) ;
assign n98 =  ( n27 ) ? ( LB2D_shift_0 ) : ( n97 ) ;
assign n99 =  ( n22 ) ? ( LB2D_shift_1 ) : ( n98 ) ;
assign n100 =  ( n13 ) ? ( LB2D_shift_0 ) : ( n99 ) ;
assign n101 =  ( n4 ) ? ( LB2D_shift_0 ) : ( n100 ) ;
assign n102 =  ( n38 ) ? ( LB2D_shift_1 ) : ( LB2D_shift_1 ) ;
assign n103 =  ( n27 ) ? ( LB2D_shift_1 ) : ( n102 ) ;
assign n104 =  ( n22 ) ? ( LB2D_shift_2 ) : ( n103 ) ;
assign n105 =  ( n13 ) ? ( LB2D_shift_1 ) : ( n104 ) ;
assign n106 =  ( n4 ) ? ( LB2D_shift_1 ) : ( n105 ) ;
assign n107 =  ( n38 ) ? ( LB2D_shift_2 ) : ( LB2D_shift_2 ) ;
assign n108 =  ( n27 ) ? ( LB2D_shift_2 ) : ( n107 ) ;
assign n109 =  ( n22 ) ? ( LB2D_shift_3 ) : ( n108 ) ;
assign n110 =  ( n13 ) ? ( LB2D_shift_2 ) : ( n109 ) ;
assign n111 =  ( n4 ) ? ( LB2D_shift_2 ) : ( n110 ) ;
assign n112 =  ( n38 ) ? ( LB2D_shift_3 ) : ( LB2D_shift_3 ) ;
assign n113 =  ( n27 ) ? ( LB2D_shift_3 ) : ( n112 ) ;
assign n114 =  ( n22 ) ? ( LB2D_shift_4 ) : ( n113 ) ;
assign n115 =  ( n13 ) ? ( LB2D_shift_3 ) : ( n114 ) ;
assign n116 =  ( n4 ) ? ( LB2D_shift_3 ) : ( n115 ) ;
assign n117 =  ( n38 ) ? ( LB2D_shift_4 ) : ( LB2D_shift_4 ) ;
assign n118 =  ( n27 ) ? ( LB2D_shift_4 ) : ( n117 ) ;
assign n119 =  ( n22 ) ? ( LB2D_shift_5 ) : ( n118 ) ;
assign n120 =  ( n13 ) ? ( LB2D_shift_4 ) : ( n119 ) ;
assign n121 =  ( n4 ) ? ( LB2D_shift_4 ) : ( n120 ) ;
assign n122 =  ( n38 ) ? ( LB2D_shift_5 ) : ( LB2D_shift_5 ) ;
assign n123 =  ( n27 ) ? ( LB2D_shift_5 ) : ( n122 ) ;
assign n124 =  ( n22 ) ? ( LB2D_shift_6 ) : ( n123 ) ;
assign n125 =  ( n13 ) ? ( LB2D_shift_5 ) : ( n124 ) ;
assign n126 =  ( n4 ) ? ( LB2D_shift_5 ) : ( n125 ) ;
assign n127 =  ( n38 ) ? ( LB2D_shift_6 ) : ( LB2D_shift_6 ) ;
assign n128 =  ( n27 ) ? ( LB2D_shift_6 ) : ( n127 ) ;
assign n129 =  ( n22 ) ? ( LB2D_shift_7 ) : ( n128 ) ;
assign n130 =  ( n13 ) ? ( LB2D_shift_6 ) : ( n129 ) ;
assign n131 =  ( n4 ) ? ( LB2D_shift_6 ) : ( n130 ) ;
assign n132 =  ( slice_stream_full ) == ( 1'd1 )  ;
assign n133 =  ( n132 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n134 =  ( n38 ) ? ( LB2D_shift_7 ) : ( LB2D_shift_7 ) ;
assign n135 =  ( n27 ) ? ( LB2D_shift_7 ) : ( n134 ) ;
assign n136 =  ( n22 ) ? ( n133 ) : ( n135 ) ;
assign n137 =  ( n13 ) ? ( LB2D_shift_7 ) : ( n136 ) ;
assign n138 =  ( n4 ) ? ( LB2D_shift_7 ) : ( n137 ) ;
assign n139 =  ( LB2D_shift_x ) == ( 9'd488 )  ;
assign n140 =  ( n14 ) & ( n139 )  ;
assign n141 =  ( n17 ) | ( n18 )  ;
assign n142 =  ( n140 ) & ( n141 )  ;
assign n143 =  ( LB2D_shift_x ) + ( 9'd1 )  ;
assign n144 =  ( n38 ) ? ( LB2D_shift_x ) : ( LB2D_shift_x ) ;
assign n145 =  ( n27 ) ? ( LB2D_shift_x ) : ( n144 ) ;
assign n146 =  ( n22 ) ? ( n143 ) : ( n145 ) ;
assign n147 =  ( n142 ) ? ( 9'd0 ) : ( n146 ) ;
assign n148 =  ( n13 ) ? ( LB2D_shift_x ) : ( n147 ) ;
assign n149 =  ( n4 ) ? ( LB2D_shift_x ) : ( n148 ) ;
assign n150 =  ( LB2D_shift_y ) < ( 10'd640 )  ;
assign n151 =  ( LB2D_shift_x ) < ( 9'd488 )  ;
assign n152 =  ( LB2D_shift_y ) + ( 10'd1 )  ;
assign n153 =  ( n151 ) ? ( LB2D_shift_y ) : ( n152 ) ;
assign n154 =  ( n150 ) ? ( n153 ) : ( 10'd640 ) ;
assign n155 =  ( n38 ) ? ( LB2D_shift_y ) : ( LB2D_shift_y ) ;
assign n156 =  ( n27 ) ? ( LB2D_shift_y ) : ( n155 ) ;
assign n157 =  ( n22 ) ? ( n154 ) : ( n156 ) ;
assign n158 =  ( n13 ) ? ( LB2D_shift_y ) : ( n157 ) ;
assign n159 =  ( n4 ) ? ( LB2D_shift_y ) : ( n158 ) ;
assign n160 =  ( stencil_stream_full ) == ( 1'd1 )  ;
assign n161 =  ( n160 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_0 ) ;
assign n162 = gb_fun(n161) ;
assign n163 =  ( n38 ) ? ( arg_0_TDATA ) : ( arg_0_TDATA ) ;
assign n164 =  ( n33 ) ? ( arg_0_TDATA ) : ( n163 ) ;
assign n165 =  ( n27 ) ? ( arg_0_TDATA ) : ( n164 ) ;
assign n166 =  ( n22 ) ? ( arg_0_TDATA ) : ( n165 ) ;
assign n167 =  ( n13 ) ? ( n162 ) : ( n166 ) ;
assign n168 =  ( n4 ) ? ( arg_0_TDATA ) : ( n167 ) ;
assign n169 =  ( gb_pp_it_8 ) == ( 1'd1 )  ;
assign n170 =  ( n169 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n171 =  ( n38 ) ? ( arg_0_TVALID ) : ( arg_0_TVALID ) ;
assign n172 =  ( n33 ) ? ( arg_0_TVALID ) : ( n171 ) ;
assign n173 =  ( n27 ) ? ( arg_0_TVALID ) : ( n172 ) ;
assign n174 =  ( n22 ) ? ( arg_0_TVALID ) : ( n173 ) ;
assign n175 =  ( n13 ) ? ( n170 ) : ( n174 ) ;
assign n176 =  ( n4 ) ? ( arg_0_TVALID ) : ( n175 ) ;
assign n177 =  ( n38 ) ? ( 1'd1 ) : ( arg_1_TREADY ) ;
assign n178 =  ( n37 ) ? ( 1'd1 ) : ( n177 ) ;
assign n179 =  ( n33 ) ? ( 1'd1 ) : ( n178 ) ;
assign n180 =  ( n27 ) ? ( arg_1_TREADY ) : ( n179 ) ;
assign n181 =  ( n22 ) ? ( arg_1_TREADY ) : ( n180 ) ;
assign n182 =  ( n13 ) ? ( arg_1_TREADY ) : ( n181 ) ;
assign n183 =  ( n4 ) ? ( 1'd0 ) : ( n182 ) ;
assign n184 =  ( gb_p_cnt ) + ( 19'd1 )  ;
assign n185 =  ( n184 ) == ( 19'd307200 )  ;
assign n186 =  ( n185 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n187 =  ( n38 ) ? ( gb_exit_it_1 ) : ( gb_exit_it_1 ) ;
assign n188 =  ( n27 ) ? ( gb_exit_it_1 ) : ( n187 ) ;
assign n189 =  ( n22 ) ? ( gb_exit_it_1 ) : ( n188 ) ;
assign n190 =  ( n13 ) ? ( n186 ) : ( n189 ) ;
assign n191 =  ( n4 ) ? ( gb_exit_it_1 ) : ( n190 ) ;
assign n192 =  ( n38 ) ? ( gb_exit_it_2 ) : ( gb_exit_it_2 ) ;
assign n193 =  ( n27 ) ? ( gb_exit_it_2 ) : ( n192 ) ;
assign n194 =  ( n22 ) ? ( gb_exit_it_2 ) : ( n193 ) ;
assign n195 =  ( n13 ) ? ( gb_exit_it_1 ) : ( n194 ) ;
assign n196 =  ( n4 ) ? ( gb_exit_it_2 ) : ( n195 ) ;
assign n197 =  ( n38 ) ? ( gb_exit_it_3 ) : ( gb_exit_it_3 ) ;
assign n198 =  ( n27 ) ? ( gb_exit_it_3 ) : ( n197 ) ;
assign n199 =  ( n22 ) ? ( gb_exit_it_3 ) : ( n198 ) ;
assign n200 =  ( n13 ) ? ( gb_exit_it_2 ) : ( n199 ) ;
assign n201 =  ( n4 ) ? ( gb_exit_it_3 ) : ( n200 ) ;
assign n202 =  ( n38 ) ? ( gb_exit_it_4 ) : ( gb_exit_it_4 ) ;
assign n203 =  ( n27 ) ? ( gb_exit_it_4 ) : ( n202 ) ;
assign n204 =  ( n22 ) ? ( gb_exit_it_4 ) : ( n203 ) ;
assign n205 =  ( n13 ) ? ( gb_exit_it_3 ) : ( n204 ) ;
assign n206 =  ( n4 ) ? ( gb_exit_it_4 ) : ( n205 ) ;
assign n207 =  ( n38 ) ? ( gb_exit_it_5 ) : ( gb_exit_it_5 ) ;
assign n208 =  ( n27 ) ? ( gb_exit_it_5 ) : ( n207 ) ;
assign n209 =  ( n22 ) ? ( gb_exit_it_5 ) : ( n208 ) ;
assign n210 =  ( n13 ) ? ( gb_exit_it_4 ) : ( n209 ) ;
assign n211 =  ( n4 ) ? ( gb_exit_it_5 ) : ( n210 ) ;
assign n212 =  ( n38 ) ? ( gb_exit_it_6 ) : ( gb_exit_it_6 ) ;
assign n213 =  ( n27 ) ? ( gb_exit_it_6 ) : ( n212 ) ;
assign n214 =  ( n22 ) ? ( gb_exit_it_6 ) : ( n213 ) ;
assign n215 =  ( n13 ) ? ( gb_exit_it_5 ) : ( n214 ) ;
assign n216 =  ( n4 ) ? ( gb_exit_it_6 ) : ( n215 ) ;
assign n217 =  ( n38 ) ? ( gb_exit_it_7 ) : ( gb_exit_it_7 ) ;
assign n218 =  ( n27 ) ? ( gb_exit_it_7 ) : ( n217 ) ;
assign n219 =  ( n22 ) ? ( gb_exit_it_7 ) : ( n218 ) ;
assign n220 =  ( n13 ) ? ( gb_exit_it_6 ) : ( n219 ) ;
assign n221 =  ( n4 ) ? ( gb_exit_it_7 ) : ( n220 ) ;
assign n222 =  ( n38 ) ? ( gb_exit_it_8 ) : ( gb_exit_it_8 ) ;
assign n223 =  ( n27 ) ? ( gb_exit_it_8 ) : ( n222 ) ;
assign n224 =  ( n22 ) ? ( gb_exit_it_8 ) : ( n223 ) ;
assign n225 =  ( n13 ) ? ( gb_exit_it_7 ) : ( n224 ) ;
assign n226 =  ( n4 ) ? ( gb_exit_it_8 ) : ( n225 ) ;
assign n227 =  ( gb_p_cnt ) < ( 19'd307200 )  ;
assign n228 =  ( n227 ) ? ( n184 ) : ( 19'd307200 ) ;
assign n229 =  ( n38 ) ? ( gb_p_cnt ) : ( gb_p_cnt ) ;
assign n230 =  ( n27 ) ? ( gb_p_cnt ) : ( n229 ) ;
assign n231 =  ( n22 ) ? ( gb_p_cnt ) : ( n230 ) ;
assign n232 =  ( n13 ) ? ( n228 ) : ( n231 ) ;
assign n233 =  ( n4 ) ? ( gb_p_cnt ) : ( n232 ) ;
assign n234 =  ( n38 ) ? ( gb_pp_it_1 ) : ( gb_pp_it_1 ) ;
assign n235 =  ( n27 ) ? ( gb_pp_it_1 ) : ( n234 ) ;
assign n236 =  ( n22 ) ? ( gb_pp_it_1 ) : ( n235 ) ;
assign n237 =  ( n13 ) ? ( 1'd1 ) : ( n236 ) ;
assign n238 =  ( n4 ) ? ( gb_pp_it_1 ) : ( n237 ) ;
assign n239 =  ( n38 ) ? ( gb_pp_it_2 ) : ( gb_pp_it_2 ) ;
assign n240 =  ( n27 ) ? ( gb_pp_it_2 ) : ( n239 ) ;
assign n241 =  ( n22 ) ? ( gb_pp_it_2 ) : ( n240 ) ;
assign n242 =  ( n13 ) ? ( gb_pp_it_1 ) : ( n241 ) ;
assign n243 =  ( n4 ) ? ( gb_pp_it_2 ) : ( n242 ) ;
assign n244 =  ( n38 ) ? ( gb_pp_it_3 ) : ( gb_pp_it_3 ) ;
assign n245 =  ( n27 ) ? ( gb_pp_it_3 ) : ( n244 ) ;
assign n246 =  ( n22 ) ? ( gb_pp_it_3 ) : ( n245 ) ;
assign n247 =  ( n13 ) ? ( gb_pp_it_2 ) : ( n246 ) ;
assign n248 =  ( n4 ) ? ( gb_pp_it_3 ) : ( n247 ) ;
assign n249 =  ( n38 ) ? ( gb_pp_it_4 ) : ( gb_pp_it_4 ) ;
assign n250 =  ( n27 ) ? ( gb_pp_it_4 ) : ( n249 ) ;
assign n251 =  ( n22 ) ? ( gb_pp_it_4 ) : ( n250 ) ;
assign n252 =  ( n13 ) ? ( gb_pp_it_3 ) : ( n251 ) ;
assign n253 =  ( n4 ) ? ( gb_pp_it_4 ) : ( n252 ) ;
assign n254 =  ( n38 ) ? ( gb_pp_it_5 ) : ( gb_pp_it_5 ) ;
assign n255 =  ( n27 ) ? ( gb_pp_it_5 ) : ( n254 ) ;
assign n256 =  ( n22 ) ? ( gb_pp_it_5 ) : ( n255 ) ;
assign n257 =  ( n13 ) ? ( gb_pp_it_4 ) : ( n256 ) ;
assign n258 =  ( n4 ) ? ( gb_pp_it_5 ) : ( n257 ) ;
assign n259 =  ( n38 ) ? ( gb_pp_it_6 ) : ( gb_pp_it_6 ) ;
assign n260 =  ( n27 ) ? ( gb_pp_it_6 ) : ( n259 ) ;
assign n261 =  ( n22 ) ? ( gb_pp_it_6 ) : ( n260 ) ;
assign n262 =  ( n13 ) ? ( gb_pp_it_5 ) : ( n261 ) ;
assign n263 =  ( n4 ) ? ( gb_pp_it_6 ) : ( n262 ) ;
assign n264 =  ( n38 ) ? ( gb_pp_it_7 ) : ( gb_pp_it_7 ) ;
assign n265 =  ( n27 ) ? ( gb_pp_it_7 ) : ( n264 ) ;
assign n266 =  ( n22 ) ? ( gb_pp_it_7 ) : ( n265 ) ;
assign n267 =  ( n13 ) ? ( gb_pp_it_6 ) : ( n266 ) ;
assign n268 =  ( n4 ) ? ( gb_pp_it_7 ) : ( n267 ) ;
assign n269 =  ( n38 ) ? ( gb_pp_it_8 ) : ( gb_pp_it_8 ) ;
assign n270 =  ( n27 ) ? ( gb_pp_it_8 ) : ( n269 ) ;
assign n271 =  ( n22 ) ? ( gb_pp_it_8 ) : ( n270 ) ;
assign n272 =  ( n13 ) ? ( gb_pp_it_7 ) : ( n271 ) ;
assign n273 =  ( n4 ) ? ( gb_pp_it_8 ) : ( n272 ) ;
assign n274 =  ( n38 ) ? ( gb_pp_it_9 ) : ( gb_pp_it_9 ) ;
assign n275 =  ( n27 ) ? ( gb_pp_it_9 ) : ( n274 ) ;
assign n276 =  ( n22 ) ? ( gb_pp_it_9 ) : ( n275 ) ;
assign n277 =  ( n13 ) ? ( gb_pp_it_8 ) : ( n276 ) ;
assign n278 =  ( n4 ) ? ( gb_pp_it_9 ) : ( n277 ) ;
assign n279 =  ( n38 ) ? ( LB1D_uIn ) : ( in_stream_buff_0 ) ;
assign n280 =  ( n33 ) ? ( LB1D_uIn ) : ( n279 ) ;
assign n281 =  ( n27 ) ? ( in_stream_buff_0 ) : ( n280 ) ;
assign n282 =  ( n22 ) ? ( in_stream_buff_0 ) : ( n281 ) ;
assign n283 =  ( n13 ) ? ( in_stream_buff_0 ) : ( n282 ) ;
assign n284 =  ( n4 ) ? ( in_stream_buff_0 ) : ( n283 ) ;
assign n285 =  ( n38 ) ? ( in_stream_buff_0 ) : ( in_stream_buff_1 ) ;
assign n286 =  ( n33 ) ? ( in_stream_buff_0 ) : ( n285 ) ;
assign n287 =  ( n27 ) ? ( in_stream_buff_1 ) : ( n286 ) ;
assign n288 =  ( n22 ) ? ( in_stream_buff_1 ) : ( n287 ) ;
assign n289 =  ( n13 ) ? ( in_stream_buff_1 ) : ( n288 ) ;
assign n290 =  ( n4 ) ? ( in_stream_buff_1 ) : ( n289 ) ;
assign n291 =  ( in_stream_full ) == ( 1'd1 )  ;
assign n292 =  ( n291 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n293 =  ( n38 ) ? ( 1'd0 ) : ( in_stream_empty ) ;
assign n294 =  ( n33 ) ? ( 1'd0 ) : ( n293 ) ;
assign n295 =  ( n27 ) ? ( n292 ) : ( n294 ) ;
assign n296 =  ( n22 ) ? ( in_stream_empty ) : ( n295 ) ;
assign n297 =  ( n13 ) ? ( in_stream_empty ) : ( n296 ) ;
assign n298 =  ( n4 ) ? ( in_stream_empty ) : ( n297 ) ;
assign n299 =  ( in_stream_empty ) == ( 1'd1 )  ;
assign n300 =  ( n299 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n301 =  ( n38 ) ? ( n300 ) : ( in_stream_full ) ;
assign n302 =  ( n33 ) ? ( n300 ) : ( n301 ) ;
assign n303 =  ( n27 ) ? ( 1'd0 ) : ( n302 ) ;
assign n304 =  ( n22 ) ? ( in_stream_full ) : ( n303 ) ;
assign n305 =  ( n13 ) ? ( in_stream_full ) : ( n304 ) ;
assign n306 =  ( n4 ) ? ( in_stream_full ) : ( n305 ) ;
assign n307 =  ( n291 ) ? ( in_stream_buff_1 ) : ( in_stream_buff_0 ) ;
assign n308 =  ( LB2D_proc_w ) == ( 64'd0 )  ;
assign n309 =  ( LB2D_proc_x ) - ( 9'd1 )  ;
assign n310 =  (  LB2D_proc_7 [ n309 ] )  ;
assign n311 =  ( LB2D_proc_w ) == ( 64'd1 )  ;
assign n312 =  (  LB2D_proc_0 [ n309 ] )  ;
assign n313 =  ( LB2D_proc_w ) == ( 64'd2 )  ;
assign n314 =  (  LB2D_proc_1 [ n309 ] )  ;
assign n315 =  ( LB2D_proc_w ) == ( 64'd3 )  ;
assign n316 =  (  LB2D_proc_2 [ n309 ] )  ;
assign n317 =  ( LB2D_proc_w ) == ( 64'd4 )  ;
assign n318 =  (  LB2D_proc_3 [ n309 ] )  ;
assign n319 =  ( LB2D_proc_w ) == ( 64'd5 )  ;
assign n320 =  (  LB2D_proc_4 [ n309 ] )  ;
assign n321 =  ( LB2D_proc_w ) == ( 64'd6 )  ;
assign n322 =  (  LB2D_proc_5 [ n309 ] )  ;
assign n323 =  (  LB2D_proc_6 [ n309 ] )  ;
assign n324 =  ( n321 ) ? ( n322 ) : ( n323 ) ;
assign n325 =  ( n319 ) ? ( n320 ) : ( n324 ) ;
assign n326 =  ( n317 ) ? ( n318 ) : ( n325 ) ;
assign n327 =  ( n315 ) ? ( n316 ) : ( n326 ) ;
assign n328 =  ( n313 ) ? ( n314 ) : ( n327 ) ;
assign n329 =  ( n311 ) ? ( n312 ) : ( n328 ) ;
assign n330 =  ( n308 ) ? ( n310 ) : ( n329 ) ;
assign n331 =  ( n321 ) ? ( n320 ) : ( n322 ) ;
assign n332 =  ( n319 ) ? ( n318 ) : ( n331 ) ;
assign n333 =  ( n317 ) ? ( n316 ) : ( n332 ) ;
assign n334 =  ( n315 ) ? ( n314 ) : ( n333 ) ;
assign n335 =  ( n313 ) ? ( n312 ) : ( n334 ) ;
assign n336 =  ( n311 ) ? ( n310 ) : ( n335 ) ;
assign n337 =  ( n308 ) ? ( n323 ) : ( n336 ) ;
assign n338 =  ( n321 ) ? ( n318 ) : ( n320 ) ;
assign n339 =  ( n319 ) ? ( n316 ) : ( n338 ) ;
assign n340 =  ( n317 ) ? ( n314 ) : ( n339 ) ;
assign n341 =  ( n315 ) ? ( n312 ) : ( n340 ) ;
assign n342 =  ( n313 ) ? ( n310 ) : ( n341 ) ;
assign n343 =  ( n311 ) ? ( n323 ) : ( n342 ) ;
assign n344 =  ( n308 ) ? ( n322 ) : ( n343 ) ;
assign n345 =  ( n321 ) ? ( n316 ) : ( n318 ) ;
assign n346 =  ( n319 ) ? ( n314 ) : ( n345 ) ;
assign n347 =  ( n317 ) ? ( n312 ) : ( n346 ) ;
assign n348 =  ( n315 ) ? ( n310 ) : ( n347 ) ;
assign n349 =  ( n313 ) ? ( n323 ) : ( n348 ) ;
assign n350 =  ( n311 ) ? ( n322 ) : ( n349 ) ;
assign n351 =  ( n308 ) ? ( n320 ) : ( n350 ) ;
assign n352 =  ( n321 ) ? ( n314 ) : ( n316 ) ;
assign n353 =  ( n319 ) ? ( n312 ) : ( n352 ) ;
assign n354 =  ( n317 ) ? ( n310 ) : ( n353 ) ;
assign n355 =  ( n315 ) ? ( n323 ) : ( n354 ) ;
assign n356 =  ( n313 ) ? ( n322 ) : ( n355 ) ;
assign n357 =  ( n311 ) ? ( n320 ) : ( n356 ) ;
assign n358 =  ( n308 ) ? ( n318 ) : ( n357 ) ;
assign n359 =  ( n321 ) ? ( n312 ) : ( n314 ) ;
assign n360 =  ( n319 ) ? ( n310 ) : ( n359 ) ;
assign n361 =  ( n317 ) ? ( n323 ) : ( n360 ) ;
assign n362 =  ( n315 ) ? ( n322 ) : ( n361 ) ;
assign n363 =  ( n313 ) ? ( n320 ) : ( n362 ) ;
assign n364 =  ( n311 ) ? ( n318 ) : ( n363 ) ;
assign n365 =  ( n308 ) ? ( n316 ) : ( n364 ) ;
assign n366 =  ( n321 ) ? ( n310 ) : ( n312 ) ;
assign n367 =  ( n319 ) ? ( n323 ) : ( n366 ) ;
assign n368 =  ( n317 ) ? ( n322 ) : ( n367 ) ;
assign n369 =  ( n315 ) ? ( n320 ) : ( n368 ) ;
assign n370 =  ( n313 ) ? ( n318 ) : ( n369 ) ;
assign n371 =  ( n311 ) ? ( n316 ) : ( n370 ) ;
assign n372 =  ( n308 ) ? ( n314 ) : ( n371 ) ;
assign n373 =  ( n321 ) ? ( n323 ) : ( n310 ) ;
assign n374 =  ( n319 ) ? ( n322 ) : ( n373 ) ;
assign n375 =  ( n317 ) ? ( n320 ) : ( n374 ) ;
assign n376 =  ( n315 ) ? ( n318 ) : ( n375 ) ;
assign n377 =  ( n313 ) ? ( n316 ) : ( n376 ) ;
assign n378 =  ( n311 ) ? ( n314 ) : ( n377 ) ;
assign n379 =  ( n308 ) ? ( n312 ) : ( n378 ) ;
assign n380 =  { ( n372 ) , ( n379 ) }  ;
assign n381 =  { ( n365 ) , ( n380 ) }  ;
assign n382 =  { ( n358 ) , ( n381 ) }  ;
assign n383 =  { ( n351 ) , ( n382 ) }  ;
assign n384 =  { ( n344 ) , ( n383 ) }  ;
assign n385 =  { ( n337 ) , ( n384 ) }  ;
assign n386 =  { ( n330 ) , ( n385 ) }  ;
assign n387 =  { ( n307 ) , ( n386 ) }  ;
assign n388 =  ( n25 ) ? ( slice_stream_buff_0 ) : ( n387 ) ;
assign n389 =  ( n38 ) ? ( slice_stream_buff_0 ) : ( slice_stream_buff_0 ) ;
assign n390 =  ( n27 ) ? ( n388 ) : ( n389 ) ;
assign n391 =  ( n22 ) ? ( slice_stream_buff_0 ) : ( n390 ) ;
assign n392 =  ( n13 ) ? ( slice_stream_buff_0 ) : ( n391 ) ;
assign n393 =  ( n4 ) ? ( slice_stream_buff_0 ) : ( n392 ) ;
assign n394 =  ( n25 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n395 =  ( n38 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_1 ) ;
assign n396 =  ( n27 ) ? ( n394 ) : ( n395 ) ;
assign n397 =  ( n22 ) ? ( slice_stream_buff_1 ) : ( n396 ) ;
assign n398 =  ( n13 ) ? ( slice_stream_buff_1 ) : ( n397 ) ;
assign n399 =  ( n4 ) ? ( slice_stream_buff_1 ) : ( n398 ) ;
assign n400 =  ( n132 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n401 =  ( n25 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n402 =  ( n38 ) ? ( slice_stream_empty ) : ( slice_stream_empty ) ;
assign n403 =  ( n27 ) ? ( n401 ) : ( n402 ) ;
assign n404 =  ( n22 ) ? ( n400 ) : ( n403 ) ;
assign n405 =  ( n13 ) ? ( slice_stream_empty ) : ( n404 ) ;
assign n406 =  ( n4 ) ? ( slice_stream_empty ) : ( n405 ) ;
assign n407 =  ( slice_stream_empty ) == ( 1'd1 )  ;
assign n408 =  ( n407 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n409 =  ( n25 ) ? ( 1'd0 ) : ( n408 ) ;
assign n410 =  ( n38 ) ? ( slice_stream_full ) : ( slice_stream_full ) ;
assign n411 =  ( n27 ) ? ( n409 ) : ( n410 ) ;
assign n412 =  ( n22 ) ? ( 1'd0 ) : ( n411 ) ;
assign n413 =  ( n13 ) ? ( slice_stream_full ) : ( n412 ) ;
assign n414 =  ( n4 ) ? ( slice_stream_full ) : ( n413 ) ;
assign n415 =  ( LB2D_shift_x ) >= ( 9'd8 )  ;
assign n416 =  ( LB2D_shift_x ) == ( 9'd0 )  ;
assign n417 =  ( n415 ) | ( n416 )  ;
assign n418 = n133[71:64] ;
assign n419 = LB2D_shift_7[71:64] ;
assign n420 = LB2D_shift_6[71:64] ;
assign n421 = LB2D_shift_5[71:64] ;
assign n422 = LB2D_shift_4[71:64] ;
assign n423 = LB2D_shift_3[71:64] ;
assign n424 = LB2D_shift_2[71:64] ;
assign n425 = LB2D_shift_1[71:64] ;
assign n426 = LB2D_shift_0[71:64] ;
assign n427 =  { ( n425 ) , ( n426 ) }  ;
assign n428 =  { ( n424 ) , ( n427 ) }  ;
assign n429 =  { ( n423 ) , ( n428 ) }  ;
assign n430 =  { ( n422 ) , ( n429 ) }  ;
assign n431 =  { ( n421 ) , ( n430 ) }  ;
assign n432 =  { ( n420 ) , ( n431 ) }  ;
assign n433 =  { ( n419 ) , ( n432 ) }  ;
assign n434 =  { ( n418 ) , ( n433 ) }  ;
assign n435 = n133[63:56] ;
assign n436 = LB2D_shift_7[63:56] ;
assign n437 = LB2D_shift_6[63:56] ;
assign n438 = LB2D_shift_5[63:56] ;
assign n439 = LB2D_shift_4[63:56] ;
assign n440 = LB2D_shift_3[63:56] ;
assign n441 = LB2D_shift_2[63:56] ;
assign n442 = LB2D_shift_1[63:56] ;
assign n443 = LB2D_shift_0[63:56] ;
assign n444 =  { ( n442 ) , ( n443 ) }  ;
assign n445 =  { ( n441 ) , ( n444 ) }  ;
assign n446 =  { ( n440 ) , ( n445 ) }  ;
assign n447 =  { ( n439 ) , ( n446 ) }  ;
assign n448 =  { ( n438 ) , ( n447 ) }  ;
assign n449 =  { ( n437 ) , ( n448 ) }  ;
assign n450 =  { ( n436 ) , ( n449 ) }  ;
assign n451 =  { ( n435 ) , ( n450 ) }  ;
assign n452 = n133[55:48] ;
assign n453 = LB2D_shift_7[55:48] ;
assign n454 = LB2D_shift_6[55:48] ;
assign n455 = LB2D_shift_5[55:48] ;
assign n456 = LB2D_shift_4[55:48] ;
assign n457 = LB2D_shift_3[55:48] ;
assign n458 = LB2D_shift_2[55:48] ;
assign n459 = LB2D_shift_1[55:48] ;
assign n460 = LB2D_shift_0[55:48] ;
assign n461 =  { ( n459 ) , ( n460 ) }  ;
assign n462 =  { ( n458 ) , ( n461 ) }  ;
assign n463 =  { ( n457 ) , ( n462 ) }  ;
assign n464 =  { ( n456 ) , ( n463 ) }  ;
assign n465 =  { ( n455 ) , ( n464 ) }  ;
assign n466 =  { ( n454 ) , ( n465 ) }  ;
assign n467 =  { ( n453 ) , ( n466 ) }  ;
assign n468 =  { ( n452 ) , ( n467 ) }  ;
assign n469 = n133[47:40] ;
assign n470 = LB2D_shift_7[47:40] ;
assign n471 = LB2D_shift_6[47:40] ;
assign n472 = LB2D_shift_5[47:40] ;
assign n473 = LB2D_shift_4[47:40] ;
assign n474 = LB2D_shift_3[47:40] ;
assign n475 = LB2D_shift_2[47:40] ;
assign n476 = LB2D_shift_1[47:40] ;
assign n477 = LB2D_shift_0[47:40] ;
assign n478 =  { ( n476 ) , ( n477 ) }  ;
assign n479 =  { ( n475 ) , ( n478 ) }  ;
assign n480 =  { ( n474 ) , ( n479 ) }  ;
assign n481 =  { ( n473 ) , ( n480 ) }  ;
assign n482 =  { ( n472 ) , ( n481 ) }  ;
assign n483 =  { ( n471 ) , ( n482 ) }  ;
assign n484 =  { ( n470 ) , ( n483 ) }  ;
assign n485 =  { ( n469 ) , ( n484 ) }  ;
assign n486 = n133[39:32] ;
assign n487 = LB2D_shift_7[39:32] ;
assign n488 = LB2D_shift_6[39:32] ;
assign n489 = LB2D_shift_5[39:32] ;
assign n490 = LB2D_shift_4[39:32] ;
assign n491 = LB2D_shift_3[39:32] ;
assign n492 = LB2D_shift_2[39:32] ;
assign n493 = LB2D_shift_1[39:32] ;
assign n494 = LB2D_shift_0[39:32] ;
assign n495 =  { ( n493 ) , ( n494 ) }  ;
assign n496 =  { ( n492 ) , ( n495 ) }  ;
assign n497 =  { ( n491 ) , ( n496 ) }  ;
assign n498 =  { ( n490 ) , ( n497 ) }  ;
assign n499 =  { ( n489 ) , ( n498 ) }  ;
assign n500 =  { ( n488 ) , ( n499 ) }  ;
assign n501 =  { ( n487 ) , ( n500 ) }  ;
assign n502 =  { ( n486 ) , ( n501 ) }  ;
assign n503 = n133[31:24] ;
assign n504 = LB2D_shift_7[31:24] ;
assign n505 = LB2D_shift_6[31:24] ;
assign n506 = LB2D_shift_5[31:24] ;
assign n507 = LB2D_shift_4[31:24] ;
assign n508 = LB2D_shift_3[31:24] ;
assign n509 = LB2D_shift_2[31:24] ;
assign n510 = LB2D_shift_1[31:24] ;
assign n511 = LB2D_shift_0[31:24] ;
assign n512 =  { ( n510 ) , ( n511 ) }  ;
assign n513 =  { ( n509 ) , ( n512 ) }  ;
assign n514 =  { ( n508 ) , ( n513 ) }  ;
assign n515 =  { ( n507 ) , ( n514 ) }  ;
assign n516 =  { ( n506 ) , ( n515 ) }  ;
assign n517 =  { ( n505 ) , ( n516 ) }  ;
assign n518 =  { ( n504 ) , ( n517 ) }  ;
assign n519 =  { ( n503 ) , ( n518 ) }  ;
assign n520 = n133[23:16] ;
assign n521 = LB2D_shift_7[23:16] ;
assign n522 = LB2D_shift_6[23:16] ;
assign n523 = LB2D_shift_5[23:16] ;
assign n524 = LB2D_shift_4[23:16] ;
assign n525 = LB2D_shift_3[23:16] ;
assign n526 = LB2D_shift_2[23:16] ;
assign n527 = LB2D_shift_1[23:16] ;
assign n528 = LB2D_shift_0[23:16] ;
assign n529 =  { ( n527 ) , ( n528 ) }  ;
assign n530 =  { ( n526 ) , ( n529 ) }  ;
assign n531 =  { ( n525 ) , ( n530 ) }  ;
assign n532 =  { ( n524 ) , ( n531 ) }  ;
assign n533 =  { ( n523 ) , ( n532 ) }  ;
assign n534 =  { ( n522 ) , ( n533 ) }  ;
assign n535 =  { ( n521 ) , ( n534 ) }  ;
assign n536 =  { ( n520 ) , ( n535 ) }  ;
assign n537 = n133[15:8] ;
assign n538 = LB2D_shift_7[15:8] ;
assign n539 = LB2D_shift_6[15:8] ;
assign n540 = LB2D_shift_5[15:8] ;
assign n541 = LB2D_shift_4[15:8] ;
assign n542 = LB2D_shift_3[15:8] ;
assign n543 = LB2D_shift_2[15:8] ;
assign n544 = LB2D_shift_1[15:8] ;
assign n545 = LB2D_shift_0[15:8] ;
assign n546 =  { ( n544 ) , ( n545 ) }  ;
assign n547 =  { ( n543 ) , ( n546 ) }  ;
assign n548 =  { ( n542 ) , ( n547 ) }  ;
assign n549 =  { ( n541 ) , ( n548 ) }  ;
assign n550 =  { ( n540 ) , ( n549 ) }  ;
assign n551 =  { ( n539 ) , ( n550 ) }  ;
assign n552 =  { ( n538 ) , ( n551 ) }  ;
assign n553 =  { ( n537 ) , ( n552 ) }  ;
assign n554 = n133[7:0] ;
assign n555 = LB2D_shift_7[7:0] ;
assign n556 = LB2D_shift_6[7:0] ;
assign n557 = LB2D_shift_5[7:0] ;
assign n558 = LB2D_shift_4[7:0] ;
assign n559 = LB2D_shift_3[7:0] ;
assign n560 = LB2D_shift_2[7:0] ;
assign n561 = LB2D_shift_1[7:0] ;
assign n562 = LB2D_shift_0[7:0] ;
assign n563 =  { ( n561 ) , ( n562 ) }  ;
assign n564 =  { ( n560 ) , ( n563 ) }  ;
assign n565 =  { ( n559 ) , ( n564 ) }  ;
assign n566 =  { ( n558 ) , ( n565 ) }  ;
assign n567 =  { ( n557 ) , ( n566 ) }  ;
assign n568 =  { ( n556 ) , ( n567 ) }  ;
assign n569 =  { ( n555 ) , ( n568 ) }  ;
assign n570 =  { ( n554 ) , ( n569 ) }  ;
assign n571 =  { ( n553 ) , ( n570 ) }  ;
assign n572 =  { ( n536 ) , ( n571 ) }  ;
assign n573 =  { ( n519 ) , ( n572 ) }  ;
assign n574 =  { ( n502 ) , ( n573 ) }  ;
assign n575 =  { ( n485 ) , ( n574 ) }  ;
assign n576 =  { ( n468 ) , ( n575 ) }  ;
assign n577 =  { ( n451 ) , ( n576 ) }  ;
assign n578 =  { ( n434 ) , ( n577 ) }  ;
assign n579 =  ( n417 ) ? ( n578 ) : ( stencil_stream_buff_0 ) ;
assign n580 =  ( n38 ) ? ( stencil_stream_buff_0 ) : ( stencil_stream_buff_0 ) ;
assign n581 =  ( n27 ) ? ( stencil_stream_buff_0 ) : ( n580 ) ;
assign n582 =  ( n22 ) ? ( n579 ) : ( n581 ) ;
assign n583 =  ( n13 ) ? ( stencil_stream_buff_0 ) : ( n582 ) ;
assign n584 =  ( n4 ) ? ( stencil_stream_buff_0 ) : ( n583 ) ;
assign n585 =  ( n38 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_1 ) ;
assign n586 =  ( n27 ) ? ( stencil_stream_buff_1 ) : ( n585 ) ;
assign n587 =  ( n22 ) ? ( stencil_stream_buff_0 ) : ( n586 ) ;
assign n588 =  ( n13 ) ? ( stencil_stream_buff_1 ) : ( n587 ) ;
assign n589 =  ( n4 ) ? ( stencil_stream_buff_1 ) : ( n588 ) ;
assign n590 =  ( n160 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n591 = ~ ( n417 ) ;
assign n592 =  ( n591 ) ? ( stencil_stream_empty ) : ( 1'd0 ) ;
assign n593 =  ( n38 ) ? ( stencil_stream_empty ) : ( stencil_stream_empty ) ;
assign n594 =  ( n27 ) ? ( stencil_stream_empty ) : ( n593 ) ;
assign n595 =  ( n22 ) ? ( n592 ) : ( n594 ) ;
assign n596 =  ( n13 ) ? ( n590 ) : ( n595 ) ;
assign n597 =  ( n4 ) ? ( stencil_stream_empty ) : ( n596 ) ;
assign n598 =  ( n9 ) ? ( 1'd0 ) : ( 1'd0 ) ;
assign n599 =  ( stencil_stream_empty ) == ( 1'd1 )  ;
assign n600 =  ( n599 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n601 =  ( n591 ) ? ( stencil_stream_full ) : ( n600 ) ;
assign n602 =  ( n38 ) ? ( stencil_stream_full ) : ( stencil_stream_full ) ;
assign n603 =  ( n27 ) ? ( stencil_stream_full ) : ( n602 ) ;
assign n604 =  ( n22 ) ? ( n601 ) : ( n603 ) ;
assign n605 =  ( n13 ) ? ( n598 ) : ( n604 ) ;
assign n606 =  ( n4 ) ? ( stencil_stream_full ) : ( n605 ) ;
assign n607 = ~ ( n4 ) ;
assign n608 = ~ ( n13 ) ;
assign n609 =  ( n607 ) & ( n608 )  ;
assign n610 = ~ ( n22 ) ;
assign n611 =  ( n609 ) & ( n610 )  ;
assign n612 = ~ ( n27 ) ;
assign n613 =  ( n611 ) & ( n612 )  ;
assign n614 = ~ ( n38 ) ;
assign n615 =  ( n613 ) & ( n614 )  ;
assign n616 =  ( n613 ) & ( n38 )  ;
assign n617 =  ( n611 ) & ( n27 )  ;
assign n618 = ~ ( n308 ) ;
assign n619 =  ( n617 ) & ( n618 )  ;
assign n620 =  ( n617 ) & ( n308 )  ;
assign n621 =  ( n609 ) & ( n22 )  ;
assign n622 =  ( n607 ) & ( n13 )  ;
assign LB2D_proc_0_addr0 = n620 ? (n309) : (0);
assign LB2D_proc_0_data0 = n620 ? (n307) : (LB2D_proc_0[0]);
assign n623 = ~ ( n311 ) ;
assign n624 =  ( n617 ) & ( n623 )  ;
assign n625 =  ( n617 ) & ( n311 )  ;
assign LB2D_proc_1_addr0 = n625 ? (n309) : (0);
assign LB2D_proc_1_data0 = n625 ? (n307) : (LB2D_proc_1[0]);
assign n626 = ~ ( n313 ) ;
assign n627 =  ( n617 ) & ( n626 )  ;
assign n628 =  ( n617 ) & ( n313 )  ;
assign LB2D_proc_2_addr0 = n628 ? (n309) : (0);
assign LB2D_proc_2_data0 = n628 ? (n307) : (LB2D_proc_2[0]);
assign n629 = ~ ( n315 ) ;
assign n630 =  ( n617 ) & ( n629 )  ;
assign n631 =  ( n617 ) & ( n315 )  ;
assign LB2D_proc_3_addr0 = n631 ? (n309) : (0);
assign LB2D_proc_3_data0 = n631 ? (n307) : (LB2D_proc_3[0]);
assign n632 = ~ ( n317 ) ;
assign n633 =  ( n617 ) & ( n632 )  ;
assign n634 =  ( n617 ) & ( n317 )  ;
assign LB2D_proc_4_addr0 = n634 ? (n309) : (0);
assign LB2D_proc_4_data0 = n634 ? (n307) : (LB2D_proc_4[0]);
assign n635 = ~ ( n319 ) ;
assign n636 =  ( n617 ) & ( n635 )  ;
assign n637 =  ( n617 ) & ( n319 )  ;
assign LB2D_proc_5_addr0 = n637 ? (n309) : (0);
assign LB2D_proc_5_data0 = n637 ? (n307) : (LB2D_proc_5[0]);
assign n638 = ~ ( n321 ) ;
assign n639 =  ( n617 ) & ( n638 )  ;
assign n640 =  ( n617 ) & ( n321 )  ;
assign LB2D_proc_6_addr0 = n640 ? (n309) : (0);
assign LB2D_proc_6_data0 = n640 ? (n307) : (LB2D_proc_6[0]);
assign n641 = ~ ( n72 ) ;
assign n642 =  ( n617 ) & ( n641 )  ;
assign n643 =  ( n617 ) & ( n72 )  ;
assign LB2D_proc_7_addr0 = n643 ? (n309) : (0);
assign LB2D_proc_7_data0 = n643 ? (n307) : (LB2D_proc_7[0]);
/*
function [7:0] gb_fun ;
input [647:0] arg0;
    begin
//TODO: Add the specific function HERE.    end
endfunction
*/

always @(posedge clk) begin
   if(rst) begin
       LB1D_buff <= LB1D_buff;
       LB1D_in <= LB1D_in;
       LB1D_it_1 <= LB1D_it_1;
       LB1D_p_cnt <= LB1D_p_cnt;
       LB1D_uIn <= LB1D_uIn;
       LB2D_proc_w <= LB2D_proc_w;
       LB2D_proc_x <= LB2D_proc_x;
       LB2D_proc_y <= LB2D_proc_y;
       LB2D_shift_0 <= LB2D_shift_0;
       LB2D_shift_1 <= LB2D_shift_1;
       LB2D_shift_2 <= LB2D_shift_2;
       LB2D_shift_3 <= LB2D_shift_3;
       LB2D_shift_4 <= LB2D_shift_4;
       LB2D_shift_5 <= LB2D_shift_5;
       LB2D_shift_6 <= LB2D_shift_6;
       LB2D_shift_7 <= LB2D_shift_7;
       LB2D_shift_x <= LB2D_shift_x;
       LB2D_shift_y <= LB2D_shift_y;
       arg_0_TDATA <= arg_0_TDATA;
       arg_0_TVALID <= arg_0_TVALID;
       arg_1_TREADY <= arg_1_TREADY;
       gb_exit_it_1 <= gb_exit_it_1;
       gb_exit_it_2 <= gb_exit_it_2;
       gb_exit_it_3 <= gb_exit_it_3;
       gb_exit_it_4 <= gb_exit_it_4;
       gb_exit_it_5 <= gb_exit_it_5;
       gb_exit_it_6 <= gb_exit_it_6;
       gb_exit_it_7 <= gb_exit_it_7;
       gb_exit_it_8 <= gb_exit_it_8;
       gb_p_cnt <= gb_p_cnt;
       gb_pp_it_1 <= gb_pp_it_1;
       gb_pp_it_2 <= gb_pp_it_2;
       gb_pp_it_3 <= gb_pp_it_3;
       gb_pp_it_4 <= gb_pp_it_4;
       gb_pp_it_5 <= gb_pp_it_5;
       gb_pp_it_6 <= gb_pp_it_6;
       gb_pp_it_7 <= gb_pp_it_7;
       gb_pp_it_8 <= gb_pp_it_8;
       gb_pp_it_9 <= gb_pp_it_9;
       in_stream_buff_0 <= in_stream_buff_0;
       in_stream_buff_1 <= in_stream_buff_1;
       in_stream_empty <= in_stream_empty;
       in_stream_full <= in_stream_full;
       slice_stream_buff_0 <= slice_stream_buff_0;
       slice_stream_buff_1 <= slice_stream_buff_1;
       slice_stream_empty <= slice_stream_empty;
       slice_stream_full <= slice_stream_full;
       stencil_stream_buff_0 <= stencil_stream_buff_0;
       stencil_stream_buff_1 <= stencil_stream_buff_1;
       stencil_stream_empty <= stencil_stream_empty;
       stencil_stream_full <= stencil_stream_full;
   end
   else if(step) begin
       LB1D_buff <= n45;
       LB1D_in <= n52;
       LB1D_it_1 <= n55;
       LB1D_p_cnt <= n63;
       LB1D_uIn <= n70;
       LB2D_proc_w <= n80;
       LB2D_proc_x <= n87;
       LB2D_proc_y <= n96;
       LB2D_shift_0 <= n101;
       LB2D_shift_1 <= n106;
       LB2D_shift_2 <= n111;
       LB2D_shift_3 <= n116;
       LB2D_shift_4 <= n121;
       LB2D_shift_5 <= n126;
       LB2D_shift_6 <= n131;
       LB2D_shift_7 <= n138;
       LB2D_shift_x <= n149;
       LB2D_shift_y <= n159;
       arg_0_TDATA <= n168;
       arg_0_TVALID <= n176;
       arg_1_TREADY <= n183;
       gb_exit_it_1 <= n191;
       gb_exit_it_2 <= n196;
       gb_exit_it_3 <= n201;
       gb_exit_it_4 <= n206;
       gb_exit_it_5 <= n211;
       gb_exit_it_6 <= n216;
       gb_exit_it_7 <= n221;
       gb_exit_it_8 <= n226;
       gb_p_cnt <= n233;
       gb_pp_it_1 <= n238;
       gb_pp_it_2 <= n243;
       gb_pp_it_3 <= n248;
       gb_pp_it_4 <= n253;
       gb_pp_it_5 <= n258;
       gb_pp_it_6 <= n263;
       gb_pp_it_7 <= n268;
       gb_pp_it_8 <= n273;
       gb_pp_it_9 <= n278;
       in_stream_buff_0 <= n284;
       in_stream_buff_1 <= n290;
       in_stream_empty <= n298;
       in_stream_full <= n306;
       slice_stream_buff_0 <= n393;
       slice_stream_buff_1 <= n399;
       slice_stream_empty <= n406;
       slice_stream_full <= n414;
       stencil_stream_buff_0 <= n584;
       stencil_stream_buff_1 <= n589;
       stencil_stream_empty <= n597;
       stencil_stream_full <= n606;
       LB2D_proc_0 [ LB2D_proc_0_addr0 ] <= LB2D_proc_0_data0;
       LB2D_proc_1 [ LB2D_proc_1_addr0 ] <= LB2D_proc_1_data0;
       LB2D_proc_2 [ LB2D_proc_2_addr0 ] <= LB2D_proc_2_data0;
       LB2D_proc_3 [ LB2D_proc_3_addr0 ] <= LB2D_proc_3_data0;
       LB2D_proc_4 [ LB2D_proc_4_addr0 ] <= LB2D_proc_4_data0;
       LB2D_proc_5 [ LB2D_proc_5_addr0 ] <= LB2D_proc_5_data0;
       LB2D_proc_6 [ LB2D_proc_6_addr0 ] <= LB2D_proc_6_data0;
       LB2D_proc_7 [ LB2D_proc_7_addr0 ] <= LB2D_proc_7_data0;
   end
end
endmodule
