module GB(
arg_0_TREADY,
arg_1_TDATA,
arg_1_TVALID,
LB1D_buff,
LB1D_in,
LB1D_it_1,
LB1D_p_cnt,
LB1D_uIn,
LB2D_proc_w,
LB2D_proc_x,
LB2D_proc_y,
LB2D_shift_0,
LB2D_shift_1,
LB2D_shift_2,
LB2D_shift_3,
LB2D_shift_4,
LB2D_shift_5,
LB2D_shift_6,
LB2D_shift_7,
LB2D_shift_x,
LB2D_shift_y,
arg_0_TDATA,
arg_0_TVALID,
arg_1_TREADY,
gb_exit_it_1,
gb_exit_it_2,
gb_exit_it_3,
gb_exit_it_4,
gb_exit_it_5,
gb_exit_it_6,
gb_exit_it_7,
gb_exit_it_8,
gb_p_cnt,
gb_pp_it_1,
gb_pp_it_2,
gb_pp_it_3,
gb_pp_it_4,
gb_pp_it_5,
gb_pp_it_6,
gb_pp_it_7,
gb_pp_it_8,
gb_pp_it_9,
in_stream_buff_0,
in_stream_buff_1,
in_stream_empty,
in_stream_full,
slice_stream_buff_0,
slice_stream_buff_1,
slice_stream_empty,
slice_stream_full,
stencil_stream_buff_0,
stencil_stream_buff_1,
stencil_stream_empty,
stencil_stream_full,
clk,rst,
step
);
input            arg_0_TREADY;
input      [7:0] arg_1_TDATA;
input            arg_1_TVALID;
input clk;
input rst;
input step;
output      [7:0] LB1D_buff;
output      [7:0] LB1D_in;
output            LB1D_it_1;
output     [18:0] LB1D_p_cnt;
output      [7:0] LB1D_uIn;
output     [63:0] LB2D_proc_w;
output      [8:0] LB2D_proc_x;
output      [9:0] LB2D_proc_y;
output     [71:0] LB2D_shift_0;
output     [71:0] LB2D_shift_1;
output     [71:0] LB2D_shift_2;
output     [71:0] LB2D_shift_3;
output     [71:0] LB2D_shift_4;
output     [71:0] LB2D_shift_5;
output     [71:0] LB2D_shift_6;
output     [71:0] LB2D_shift_7;
output      [8:0] LB2D_shift_x;
output      [9:0] LB2D_shift_y;
output      [7:0] arg_0_TDATA;
output            arg_0_TVALID;
output            arg_1_TREADY;
output            gb_exit_it_1;
output            gb_exit_it_2;
output            gb_exit_it_3;
output            gb_exit_it_4;
output            gb_exit_it_5;
output            gb_exit_it_6;
output            gb_exit_it_7;
output            gb_exit_it_8;
output     [18:0] gb_p_cnt;
output            gb_pp_it_1;
output            gb_pp_it_2;
output            gb_pp_it_3;
output            gb_pp_it_4;
output            gb_pp_it_5;
output            gb_pp_it_6;
output            gb_pp_it_7;
output            gb_pp_it_8;
output            gb_pp_it_9;
output      [7:0] in_stream_buff_0;
output      [7:0] in_stream_buff_1;
output            in_stream_empty;
output            in_stream_full;
output     [71:0] slice_stream_buff_0;
output     [71:0] slice_stream_buff_1;
output            slice_stream_empty;
output            slice_stream_full;
output    [647:0] stencil_stream_buff_0;
output    [647:0] stencil_stream_buff_1;
output            stencil_stream_empty;
output            stencil_stream_full;
reg      [7:0] LB1D_buff;
reg      [7:0] LB1D_in;
reg            LB1D_it_1;
reg     [18:0] LB1D_p_cnt;
reg      [7:0] LB1D_uIn;
reg     [63:0] LB2D_proc_w;
reg      [8:0] LB2D_proc_x;
reg      [9:0] LB2D_proc_y;
reg     [71:0] LB2D_shift_0;
reg     [71:0] LB2D_shift_1;
reg     [71:0] LB2D_shift_2;
reg     [71:0] LB2D_shift_3;
reg     [71:0] LB2D_shift_4;
reg     [71:0] LB2D_shift_5;
reg     [71:0] LB2D_shift_6;
reg     [71:0] LB2D_shift_7;
reg      [8:0] LB2D_shift_x;
reg      [9:0] LB2D_shift_y;
reg      [7:0] arg_0_TDATA;
reg            arg_0_TVALID;
reg            arg_1_TREADY;
reg            gb_exit_it_1;
reg            gb_exit_it_2;
reg            gb_exit_it_3;
reg            gb_exit_it_4;
reg            gb_exit_it_5;
reg            gb_exit_it_6;
reg            gb_exit_it_7;
reg            gb_exit_it_8;
reg     [18:0] gb_p_cnt;
reg            gb_pp_it_1;
reg            gb_pp_it_2;
reg            gb_pp_it_3;
reg            gb_pp_it_4;
reg            gb_pp_it_5;
reg            gb_pp_it_6;
reg            gb_pp_it_7;
reg            gb_pp_it_8;
reg            gb_pp_it_9;
reg      [7:0] in_stream_buff_0;
reg      [7:0] in_stream_buff_1;
reg            in_stream_empty;
reg            in_stream_full;
reg     [71:0] slice_stream_buff_0;
reg     [71:0] slice_stream_buff_1;
reg            slice_stream_empty;
reg            slice_stream_full;
reg    [647:0] stencil_stream_buff_0;
reg    [647:0] stencil_stream_buff_1;
reg            stencil_stream_empty;
reg            stencil_stream_full;
wire            arg_0_TREADY;
wire      [7:0] arg_1_TDATA;
wire            arg_1_TVALID;
wire            n0;
wire            n1;
wire            n2;
wire            n3;
wire            n4;
wire            n5;
wire            n6;
wire            n7;
wire            n8;
wire            n9;
wire            n10;
wire            n11;
wire            n12;
wire            n13;
wire            n14;
wire            n15;
wire            n16;
wire            n17;
wire            n18;
wire            n19;
wire            n20;
wire            n21;
wire            n22;
wire            n23;
wire            n24;
wire            n25;
wire            n26;
wire            n27;
wire            n28;
wire            n29;
wire            n30;
wire            n31;
wire            n32;
wire            n33;
wire            n34;
wire            n35;
wire      [7:0] n36;
wire      [7:0] n37;
wire      [7:0] n38;
wire      [7:0] n39;
wire      [7:0] n40;
wire      [7:0] n41;
wire      [7:0] n42;
wire      [7:0] n43;
wire      [7:0] n44;
wire      [7:0] n45;
wire      [7:0] n46;
wire      [7:0] n47;
wire            n48;
wire            n49;
wire            n50;
wire     [18:0] n51;
wire     [18:0] n52;
wire            n53;
wire     [18:0] n54;
wire     [18:0] n55;
wire     [18:0] n56;
wire     [18:0] n57;
wire     [18:0] n58;
wire     [18:0] n59;
wire     [18:0] n60;
wire     [18:0] n61;
wire      [7:0] n62;
wire      [7:0] n63;
wire      [7:0] n64;
wire      [7:0] n65;
wire      [7:0] n66;
wire            n67;
wire            n68;
wire     [63:0] n69;
wire     [63:0] n70;
wire     [63:0] n71;
wire     [63:0] n72;
wire     [63:0] n73;
wire     [63:0] n74;
wire     [63:0] n75;
wire     [63:0] n76;
wire     [63:0] n77;
wire      [8:0] n78;
wire      [8:0] n79;
wire      [8:0] n80;
wire      [8:0] n81;
wire      [8:0] n82;
wire      [8:0] n83;
wire      [8:0] n84;
wire      [8:0] n85;
wire            n86;
wire      [9:0] n87;
wire      [9:0] n88;
wire      [9:0] n89;
wire      [9:0] n90;
wire      [9:0] n91;
wire      [9:0] n92;
wire      [9:0] n93;
wire      [9:0] n94;
wire      [9:0] n95;
wire            n96;
wire     [71:0] n97;
wire     [71:0] n98;
wire     [71:0] n99;
wire     [71:0] n100;
wire     [71:0] n101;
wire     [71:0] n102;
wire     [71:0] n103;
wire     [71:0] n104;
wire     [71:0] n105;
wire     [71:0] n106;
wire     [71:0] n107;
wire     [71:0] n108;
wire     [71:0] n109;
wire     [71:0] n110;
wire     [71:0] n111;
wire     [71:0] n112;
wire     [71:0] n113;
wire     [71:0] n114;
wire     [71:0] n115;
wire     [71:0] n116;
wire     [71:0] n117;
wire     [71:0] n118;
wire     [71:0] n119;
wire     [71:0] n120;
wire     [71:0] n121;
wire     [71:0] n122;
wire     [71:0] n123;
wire     [71:0] n124;
wire     [71:0] n125;
wire     [71:0] n126;
wire     [71:0] n127;
wire     [71:0] n128;
wire     [71:0] n129;
wire     [71:0] n130;
wire     [71:0] n131;
wire     [71:0] n132;
wire     [71:0] n133;
wire     [71:0] n134;
wire     [71:0] n135;
wire     [71:0] n136;
wire     [71:0] n137;
wire     [71:0] n138;
wire     [71:0] n139;
wire     [71:0] n140;
wire     [71:0] n141;
wire     [71:0] n142;
wire     [71:0] n143;
wire     [71:0] n144;
wire     [71:0] n145;
wire      [8:0] n146;
wire      [8:0] n147;
wire      [8:0] n148;
wire      [8:0] n149;
wire      [8:0] n150;
wire      [8:0] n151;
wire      [8:0] n152;
wire            n153;
wire            n154;
wire      [9:0] n155;
wire      [9:0] n156;
wire      [9:0] n157;
wire      [9:0] n158;
wire      [9:0] n159;
wire      [9:0] n160;
wire      [9:0] n161;
wire      [9:0] n162;
wire      [9:0] n163;
wire            n164;
wire    [647:0] n165;
wire      [7:0] n166;
wire      [7:0] n167;
wire      [7:0] n168;
wire      [7:0] n169;
wire      [7:0] n170;
wire      [7:0] n171;
wire      [7:0] n172;
wire            n173;
wire            n174;
wire            n175;
wire            n176;
wire            n177;
wire            n178;
wire            n179;
wire            n180;
wire            n181;
wire            n182;
wire            n183;
wire            n184;
wire            n185;
wire            n186;
wire            n187;
wire     [18:0] n188;
wire            n189;
wire            n190;
wire            n191;
wire            n192;
wire            n193;
wire            n194;
wire            n195;
wire            n196;
wire            n197;
wire            n198;
wire            n199;
wire            n200;
wire            n201;
wire            n202;
wire            n203;
wire            n204;
wire            n205;
wire            n206;
wire            n207;
wire            n208;
wire            n209;
wire            n210;
wire            n211;
wire            n212;
wire            n213;
wire            n214;
wire            n215;
wire            n216;
wire            n217;
wire            n218;
wire            n219;
wire            n220;
wire            n221;
wire            n222;
wire            n223;
wire            n224;
wire            n225;
wire            n226;
wire            n227;
wire            n228;
wire            n229;
wire            n230;
wire            n231;
wire            n232;
wire            n233;
wire            n234;
wire            n235;
wire            n236;
wire            n237;
wire            n238;
wire            n239;
wire     [18:0] n240;
wire     [18:0] n241;
wire     [18:0] n242;
wire     [18:0] n243;
wire     [18:0] n244;
wire     [18:0] n245;
wire     [18:0] n246;
wire            n247;
wire            n248;
wire            n249;
wire            n250;
wire            n251;
wire            n252;
wire            n253;
wire            n254;
wire            n255;
wire            n256;
wire            n257;
wire            n258;
wire            n259;
wire            n260;
wire            n261;
wire            n262;
wire            n263;
wire            n264;
wire            n265;
wire            n266;
wire            n267;
wire            n268;
wire            n269;
wire            n270;
wire            n271;
wire            n272;
wire            n273;
wire            n274;
wire            n275;
wire            n276;
wire            n277;
wire            n278;
wire            n279;
wire            n280;
wire            n281;
wire            n282;
wire            n283;
wire            n284;
wire            n285;
wire            n286;
wire            n287;
wire            n288;
wire            n289;
wire            n290;
wire            n291;
wire            n292;
wire            n293;
wire            n294;
wire            n295;
wire            n296;
wire            n297;
wire            n298;
wire            n299;
wire            n300;
wire      [7:0] n301;
wire      [7:0] n302;
wire      [7:0] n303;
wire      [7:0] n304;
wire      [7:0] n305;
wire      [7:0] n306;
wire      [7:0] n307;
wire      [7:0] n308;
wire      [7:0] n309;
wire      [7:0] n310;
wire      [7:0] n311;
wire      [7:0] n312;
wire            n313;
wire            n314;
wire            n315;
wire            n316;
wire            n317;
wire            n318;
wire            n319;
wire            n320;
wire            n321;
wire            n322;
wire            n323;
wire            n324;
wire            n325;
wire            n326;
wire            n327;
wire            n328;
wire      [7:0] n329;
wire            n330;
wire      [7:0] n331;
wire            n332;
wire      [7:0] n333;
wire            n334;
wire      [7:0] n335;
wire            n336;
wire      [7:0] n337;
wire            n338;
wire      [7:0] n339;
wire            n340;
wire      [7:0] n341;
wire            n342;
wire      [7:0] n343;
wire      [7:0] n344;
wire      [7:0] n345;
wire      [7:0] n346;
wire      [7:0] n347;
wire      [7:0] n348;
wire      [7:0] n349;
wire      [7:0] n350;
wire      [7:0] n351;
wire      [7:0] n352;
wire      [7:0] n353;
wire      [7:0] n354;
wire      [7:0] n355;
wire      [7:0] n356;
wire      [7:0] n357;
wire      [7:0] n358;
wire      [7:0] n359;
wire      [7:0] n360;
wire      [7:0] n361;
wire      [7:0] n362;
wire      [7:0] n363;
wire      [7:0] n364;
wire      [7:0] n365;
wire      [7:0] n366;
wire      [7:0] n367;
wire      [7:0] n368;
wire      [7:0] n369;
wire      [7:0] n370;
wire      [7:0] n371;
wire      [7:0] n372;
wire      [7:0] n373;
wire      [7:0] n374;
wire      [7:0] n375;
wire      [7:0] n376;
wire      [7:0] n377;
wire      [7:0] n378;
wire      [7:0] n379;
wire      [7:0] n380;
wire      [7:0] n381;
wire      [7:0] n382;
wire      [7:0] n383;
wire      [7:0] n384;
wire      [7:0] n385;
wire      [7:0] n386;
wire      [7:0] n387;
wire      [7:0] n388;
wire      [7:0] n389;
wire      [7:0] n390;
wire      [7:0] n391;
wire      [7:0] n392;
wire      [7:0] n393;
wire      [7:0] n394;
wire      [7:0] n395;
wire      [7:0] n396;
wire      [7:0] n397;
wire      [7:0] n398;
wire      [7:0] n399;
wire      [7:0] n400;
wire     [15:0] n401;
wire     [23:0] n402;
wire     [31:0] n403;
wire     [39:0] n404;
wire     [47:0] n405;
wire     [55:0] n406;
wire     [63:0] n407;
wire     [71:0] n408;
wire     [71:0] n409;
wire     [71:0] n410;
wire     [71:0] n411;
wire     [71:0] n412;
wire     [71:0] n413;
wire     [71:0] n414;
wire     [71:0] n415;
wire     [71:0] n416;
wire     [71:0] n417;
wire     [71:0] n418;
wire     [71:0] n419;
wire     [71:0] n420;
wire     [71:0] n421;
wire     [71:0] n422;
wire            n423;
wire            n424;
wire            n425;
wire            n426;
wire            n427;
wire            n428;
wire            n429;
wire            n430;
wire            n431;
wire            n432;
wire            n433;
wire            n434;
wire            n435;
wire            n436;
wire            n437;
wire            n438;
wire            n439;
wire            n440;
wire      [7:0] n441;
wire      [7:0] n442;
wire      [7:0] n443;
wire      [7:0] n444;
wire      [7:0] n445;
wire      [7:0] n446;
wire      [7:0] n447;
wire      [7:0] n448;
wire      [7:0] n449;
wire     [15:0] n450;
wire     [23:0] n451;
wire     [31:0] n452;
wire     [39:0] n453;
wire     [47:0] n454;
wire     [55:0] n455;
wire     [63:0] n456;
wire     [71:0] n457;
wire      [7:0] n458;
wire      [7:0] n459;
wire      [7:0] n460;
wire      [7:0] n461;
wire      [7:0] n462;
wire      [7:0] n463;
wire      [7:0] n464;
wire      [7:0] n465;
wire      [7:0] n466;
wire     [15:0] n467;
wire     [23:0] n468;
wire     [31:0] n469;
wire     [39:0] n470;
wire     [47:0] n471;
wire     [55:0] n472;
wire     [63:0] n473;
wire     [71:0] n474;
wire      [7:0] n475;
wire      [7:0] n476;
wire      [7:0] n477;
wire      [7:0] n478;
wire      [7:0] n479;
wire      [7:0] n480;
wire      [7:0] n481;
wire      [7:0] n482;
wire      [7:0] n483;
wire     [15:0] n484;
wire     [23:0] n485;
wire     [31:0] n486;
wire     [39:0] n487;
wire     [47:0] n488;
wire     [55:0] n489;
wire     [63:0] n490;
wire     [71:0] n491;
wire      [7:0] n492;
wire      [7:0] n493;
wire      [7:0] n494;
wire      [7:0] n495;
wire      [7:0] n496;
wire      [7:0] n497;
wire      [7:0] n498;
wire      [7:0] n499;
wire      [7:0] n500;
wire     [15:0] n501;
wire     [23:0] n502;
wire     [31:0] n503;
wire     [39:0] n504;
wire     [47:0] n505;
wire     [55:0] n506;
wire     [63:0] n507;
wire     [71:0] n508;
wire      [7:0] n509;
wire      [7:0] n510;
wire      [7:0] n511;
wire      [7:0] n512;
wire      [7:0] n513;
wire      [7:0] n514;
wire      [7:0] n515;
wire      [7:0] n516;
wire      [7:0] n517;
wire     [15:0] n518;
wire     [23:0] n519;
wire     [31:0] n520;
wire     [39:0] n521;
wire     [47:0] n522;
wire     [55:0] n523;
wire     [63:0] n524;
wire     [71:0] n525;
wire      [7:0] n526;
wire      [7:0] n527;
wire      [7:0] n528;
wire      [7:0] n529;
wire      [7:0] n530;
wire      [7:0] n531;
wire      [7:0] n532;
wire      [7:0] n533;
wire      [7:0] n534;
wire     [15:0] n535;
wire     [23:0] n536;
wire     [31:0] n537;
wire     [39:0] n538;
wire     [47:0] n539;
wire     [55:0] n540;
wire     [63:0] n541;
wire     [71:0] n542;
wire      [7:0] n543;
wire      [7:0] n544;
wire      [7:0] n545;
wire      [7:0] n546;
wire      [7:0] n547;
wire      [7:0] n548;
wire      [7:0] n549;
wire      [7:0] n550;
wire      [7:0] n551;
wire     [15:0] n552;
wire     [23:0] n553;
wire     [31:0] n554;
wire     [39:0] n555;
wire     [47:0] n556;
wire     [55:0] n557;
wire     [63:0] n558;
wire     [71:0] n559;
wire      [7:0] n560;
wire      [7:0] n561;
wire      [7:0] n562;
wire      [7:0] n563;
wire      [7:0] n564;
wire      [7:0] n565;
wire      [7:0] n566;
wire      [7:0] n567;
wire      [7:0] n568;
wire     [15:0] n569;
wire     [23:0] n570;
wire     [31:0] n571;
wire     [39:0] n572;
wire     [47:0] n573;
wire     [55:0] n574;
wire     [63:0] n575;
wire     [71:0] n576;
wire      [7:0] n577;
wire      [7:0] n578;
wire      [7:0] n579;
wire      [7:0] n580;
wire      [7:0] n581;
wire      [7:0] n582;
wire      [7:0] n583;
wire      [7:0] n584;
wire      [7:0] n585;
wire     [15:0] n586;
wire     [23:0] n587;
wire     [31:0] n588;
wire     [39:0] n589;
wire     [47:0] n590;
wire     [55:0] n591;
wire     [63:0] n592;
wire     [71:0] n593;
wire    [143:0] n594;
wire    [215:0] n595;
wire    [287:0] n596;
wire    [359:0] n597;
wire    [431:0] n598;
wire    [503:0] n599;
wire    [575:0] n600;
wire    [647:0] n601;
wire    [647:0] n602;
wire    [647:0] n603;
wire    [647:0] n604;
wire    [647:0] n605;
wire    [647:0] n606;
wire    [647:0] n607;
wire    [647:0] n608;
wire    [647:0] n609;
wire    [647:0] n610;
wire    [647:0] n611;
wire    [647:0] n612;
wire    [647:0] n613;
wire    [647:0] n614;
wire            n615;
wire            n616;
wire            n617;
wire            n618;
wire            n619;
wire            n620;
wire            n621;
wire            n622;
wire            n623;
wire            n624;
wire            n625;
wire            n626;
wire            n627;
wire            n628;
wire            n629;
wire            n630;
wire            n631;
wire            n632;
wire      [8:0] LB2D_proc_0_addr0;
wire      [7:0] LB2D_proc_0_data0;
wire            n633;
wire            n634;
wire            n635;
wire            n636;
wire            n637;
wire            n638;
wire            n639;
wire            n640;
wire            n641;
wire            n642;
wire            n643;
wire            n644;
wire            n645;
wire            n646;
wire            n647;
wire            n648;
wire            n649;
wire            n650;
wire            n651;
wire      [8:0] LB2D_proc_1_addr0;
wire      [7:0] LB2D_proc_1_data0;
wire            n652;
wire            n653;
wire            n654;
wire      [8:0] LB2D_proc_2_addr0;
wire      [7:0] LB2D_proc_2_data0;
wire            n655;
wire            n656;
wire            n657;
wire      [8:0] LB2D_proc_3_addr0;
wire      [7:0] LB2D_proc_3_data0;
wire            n658;
wire            n659;
wire            n660;
wire      [8:0] LB2D_proc_4_addr0;
wire      [7:0] LB2D_proc_4_data0;
wire            n661;
wire            n662;
wire            n663;
wire      [8:0] LB2D_proc_5_addr0;
wire      [7:0] LB2D_proc_5_data0;
wire            n664;
wire            n665;
wire            n666;
wire      [8:0] LB2D_proc_6_addr0;
wire      [7:0] LB2D_proc_6_data0;
wire            n667;
wire            n668;
wire            n669;
wire      [8:0] LB2D_proc_7_addr0;
wire      [7:0] LB2D_proc_7_data0;
wire            n670;
wire            n671;
wire            n672;
reg      [7:0] LB2D_proc_0[511:0];
reg      [7:0] LB2D_proc_1[511:0];
reg      [7:0] LB2D_proc_2[511:0];
reg      [7:0] LB2D_proc_3[511:0];
reg      [7:0] LB2D_proc_4[511:0];
reg      [7:0] LB2D_proc_5[511:0];
reg      [7:0] LB2D_proc_6[511:0];
reg      [7:0] LB2D_proc_7[511:0];
wire clk;
wire rst;
wire step;
assign n0 =  ( arg_0_TREADY ) == ( 1'd1 )  ;
assign n1 =  ( arg_0_TVALID ) == ( 1'd1 )  ;
assign n2 =  ( n0 ) & ( n1 )  ;
assign n3 =  ( arg_1_TVALID ) == ( 1'd0 )  ;
assign n4 =  ( n2 ) & ( n3 )  ;
assign n5 =  ( arg_1_TREADY ) == ( 1'd1 )  ;
assign n6 =  ( arg_1_TVALID ) == ( 1'd1 )  ;
assign n7 =  ( n5 ) & ( n6 )  ;
assign n8 =  ( arg_0_TREADY ) == ( 1'd0 )  ;
assign n9 =  ( n7 ) & ( n8 )  ;
assign n10 =  ( arg_0_TVALID ) == ( 1'd0 )  ;
assign n11 =  ( gb_exit_it_1 ) == ( 1'd0 )  ;
assign n12 =  ( stencil_stream_empty ) == ( 1'd0 )  ;
assign n13 =  ( n11 ) & ( n12 )  ;
assign n14 =  ( gb_exit_it_1 ) == ( 1'd1 )  ;
assign n15 =  ( gb_exit_it_8 ) == ( 1'd0 )  ;
assign n16 =  ( n14 ) & ( n15 )  ;
assign n17 =  ( n13 ) | ( n16 )  ;
assign n18 =  ( n10 ) & ( n17 )  ;
assign n19 =  ( slice_stream_empty ) == ( 1'd0 )  ;
assign n20 =  ( LB2D_shift_x ) != ( 9'd488 )  ;
assign n21 =  ( n19 ) & ( n20 )  ;
assign n22 =  ( stencil_stream_full ) == ( 1'd0 )  ;
assign n23 =  ( LB2D_shift_x ) < ( 9'd8 )  ;
assign n24 =  ( n22 ) | ( n23 )  ;
assign n25 =  ( n21 ) & ( n24 )  ;
assign n26 =  ( in_stream_empty ) == ( 1'd0 )  ;
assign n27 =  ( slice_stream_full ) == ( 1'd0 )  ;
assign n28 =  ( LB2D_proc_y ) < ( 10'd8 )  ;
assign n29 =  ( n27 ) | ( n28 )  ;
assign n30 =  ( n26 ) & ( n29 )  ;
assign n31 =  ( arg_1_TREADY ) == ( 1'd0 )  ;
assign n32 =  ( in_stream_full ) == ( 1'd0 )  ;
assign n33 =  ( n31 ) & ( n32 )  ;
assign n34 =  ( LB1D_it_1 ) == ( 1'd1 )  ;
assign n35 =  ( n33 ) & ( n34 )  ;
assign n36 =  ( n35 ) ? ( LB1D_uIn ) : ( LB1D_buff ) ;
assign n37 =  ( n30 ) ? ( LB1D_buff ) : ( n36 ) ;
assign n38 =  ( n25 ) ? ( LB1D_buff ) : ( n37 ) ;
assign n39 =  ( n18 ) ? ( LB1D_buff ) : ( n38 ) ;
assign n40 =  ( n9 ) ? ( LB1D_buff ) : ( n39 ) ;
assign n41 =  ( n4 ) ? ( LB1D_buff ) : ( n40 ) ;
assign n42 =  ( n35 ) ? ( LB1D_in ) : ( LB1D_in ) ;
assign n43 =  ( n30 ) ? ( LB1D_in ) : ( n42 ) ;
assign n44 =  ( n25 ) ? ( LB1D_in ) : ( n43 ) ;
assign n45 =  ( n18 ) ? ( LB1D_in ) : ( n44 ) ;
assign n46 =  ( n9 ) ? ( arg_1_TDATA ) : ( n45 ) ;
assign n47 =  ( n4 ) ? ( LB1D_in ) : ( n46 ) ;
assign n48 =  ( LB1D_it_1 ) == ( 1'd0 )  ;
assign n49 =  ( n33 ) & ( n48 )  ;
assign n50 =  ( n49 ) ? ( 1'd1 ) : ( LB1D_it_1 ) ;
assign n51 =  ( LB1D_p_cnt ) + ( 19'd1 )  ;
assign n52 =  ( 19'd316224 ) - ( 19'd1 )  ;
assign n53 =  ( LB1D_p_cnt ) == ( n52 )  ;
assign n54 =  ( n53 ) ? ( 19'd0 ) : ( n51 ) ;
assign n55 =  ( n35 ) ? ( n54 ) : ( LB1D_p_cnt ) ;
assign n56 =  ( n49 ) ? ( n51 ) : ( n55 ) ;
assign n57 =  ( n30 ) ? ( LB1D_p_cnt ) : ( n56 ) ;
assign n58 =  ( n25 ) ? ( LB1D_p_cnt ) : ( n57 ) ;
assign n59 =  ( n18 ) ? ( LB1D_p_cnt ) : ( n58 ) ;
assign n60 =  ( n9 ) ? ( LB1D_p_cnt ) : ( n59 ) ;
assign n61 =  ( n4 ) ? ( LB1D_p_cnt ) : ( n60 ) ;
assign n62 =  ( n35 ) ? ( LB1D_in ) : ( LB1D_uIn ) ;
assign n63 =  ( n30 ) ? ( LB1D_uIn ) : ( n62 ) ;
assign n64 =  ( n25 ) ? ( LB1D_uIn ) : ( n63 ) ;
assign n65 =  ( n18 ) ? ( LB1D_uIn ) : ( n64 ) ;
assign n66 =  ( n9 ) ? ( LB1D_uIn ) : ( n65 ) ;
assign n67 =  ( LB2D_proc_x ) == ( 9'd488 )  ;
assign n68 =  ( LB2D_proc_w ) == ( 64'd7 )  ;
assign n69 =  ( LB2D_proc_w ) + ( 64'd1 )  ;
assign n70 =  ( n68 ) ? ( 64'd0 ) : ( n69 ) ;
assign n71 =  ( n67 ) ? ( n70 ) : ( LB2D_proc_w ) ;
assign n72 =  ( n35 ) ? ( LB2D_proc_w ) : ( LB2D_proc_w ) ;
assign n73 =  ( n30 ) ? ( n71 ) : ( n72 ) ;
assign n74 =  ( n25 ) ? ( LB2D_proc_w ) : ( n73 ) ;
assign n75 =  ( n18 ) ? ( LB2D_proc_w ) : ( n74 ) ;
assign n76 =  ( n9 ) ? ( LB2D_proc_w ) : ( n75 ) ;
assign n77 =  ( n4 ) ? ( LB2D_proc_w ) : ( n76 ) ;
assign n78 =  ( LB2D_proc_x ) + ( 9'd1 )  ;
assign n79 =  ( n67 ) ? ( 9'd1 ) : ( n78 ) ;
assign n80 =  ( n35 ) ? ( LB2D_proc_x ) : ( LB2D_proc_x ) ;
assign n81 =  ( n30 ) ? ( n79 ) : ( n80 ) ;
assign n82 =  ( n25 ) ? ( LB2D_proc_x ) : ( n81 ) ;
assign n83 =  ( n18 ) ? ( LB2D_proc_x ) : ( n82 ) ;
assign n84 =  ( n9 ) ? ( LB2D_proc_x ) : ( n83 ) ;
assign n85 =  ( n4 ) ? ( LB2D_proc_x ) : ( n84 ) ;
assign n86 =  ( LB2D_proc_y ) == ( 10'd488 )  ;
assign n87 =  ( LB2D_proc_y ) + ( 10'd1 )  ;
assign n88 =  ( n86 ) ? ( 10'd0 ) : ( n87 ) ;
assign n89 =  ( n67 ) ? ( n88 ) : ( LB2D_proc_y ) ;
assign n90 =  ( n35 ) ? ( LB2D_proc_y ) : ( LB2D_proc_y ) ;
assign n91 =  ( n30 ) ? ( n89 ) : ( n90 ) ;
assign n92 =  ( n25 ) ? ( LB2D_proc_y ) : ( n91 ) ;
assign n93 =  ( n18 ) ? ( LB2D_proc_y ) : ( n92 ) ;
assign n94 =  ( n9 ) ? ( LB2D_proc_y ) : ( n93 ) ;
assign n95 =  ( n4 ) ? ( LB2D_proc_y ) : ( n94 ) ;
assign n96 =  ( slice_stream_full ) == ( 1'd1 )  ;
assign n97 =  ( n96 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n98 =  ( n35 ) ? ( LB2D_shift_0 ) : ( LB2D_shift_0 ) ;
assign n99 =  ( n30 ) ? ( LB2D_shift_0 ) : ( n98 ) ;
assign n100 =  ( n25 ) ? ( n97 ) : ( n99 ) ;
assign n101 =  ( n18 ) ? ( LB2D_shift_0 ) : ( n100 ) ;
assign n102 =  ( n9 ) ? ( LB2D_shift_0 ) : ( n101 ) ;
assign n103 =  ( n4 ) ? ( LB2D_shift_0 ) : ( n102 ) ;
assign n104 =  ( n35 ) ? ( LB2D_shift_1 ) : ( LB2D_shift_1 ) ;
assign n105 =  ( n30 ) ? ( LB2D_shift_1 ) : ( n104 ) ;
assign n106 =  ( n25 ) ? ( LB2D_shift_0 ) : ( n105 ) ;
assign n107 =  ( n18 ) ? ( LB2D_shift_1 ) : ( n106 ) ;
assign n108 =  ( n9 ) ? ( LB2D_shift_1 ) : ( n107 ) ;
assign n109 =  ( n4 ) ? ( LB2D_shift_1 ) : ( n108 ) ;
assign n110 =  ( n35 ) ? ( LB2D_shift_2 ) : ( LB2D_shift_2 ) ;
assign n111 =  ( n30 ) ? ( LB2D_shift_2 ) : ( n110 ) ;
assign n112 =  ( n25 ) ? ( LB2D_shift_1 ) : ( n111 ) ;
assign n113 =  ( n18 ) ? ( LB2D_shift_2 ) : ( n112 ) ;
assign n114 =  ( n9 ) ? ( LB2D_shift_2 ) : ( n113 ) ;
assign n115 =  ( n4 ) ? ( LB2D_shift_2 ) : ( n114 ) ;
assign n116 =  ( n35 ) ? ( LB2D_shift_3 ) : ( LB2D_shift_3 ) ;
assign n117 =  ( n30 ) ? ( LB2D_shift_3 ) : ( n116 ) ;
assign n118 =  ( n25 ) ? ( LB2D_shift_2 ) : ( n117 ) ;
assign n119 =  ( n18 ) ? ( LB2D_shift_3 ) : ( n118 ) ;
assign n120 =  ( n9 ) ? ( LB2D_shift_3 ) : ( n119 ) ;
assign n121 =  ( n4 ) ? ( LB2D_shift_3 ) : ( n120 ) ;
assign n122 =  ( n35 ) ? ( LB2D_shift_4 ) : ( LB2D_shift_4 ) ;
assign n123 =  ( n30 ) ? ( LB2D_shift_4 ) : ( n122 ) ;
assign n124 =  ( n25 ) ? ( LB2D_shift_3 ) : ( n123 ) ;
assign n125 =  ( n18 ) ? ( LB2D_shift_4 ) : ( n124 ) ;
assign n126 =  ( n9 ) ? ( LB2D_shift_4 ) : ( n125 ) ;
assign n127 =  ( n4 ) ? ( LB2D_shift_4 ) : ( n126 ) ;
assign n128 =  ( n35 ) ? ( LB2D_shift_5 ) : ( LB2D_shift_5 ) ;
assign n129 =  ( n30 ) ? ( LB2D_shift_5 ) : ( n128 ) ;
assign n130 =  ( n25 ) ? ( LB2D_shift_4 ) : ( n129 ) ;
assign n131 =  ( n18 ) ? ( LB2D_shift_5 ) : ( n130 ) ;
assign n132 =  ( n9 ) ? ( LB2D_shift_5 ) : ( n131 ) ;
assign n133 =  ( n4 ) ? ( LB2D_shift_5 ) : ( n132 ) ;
assign n134 =  ( n35 ) ? ( LB2D_shift_6 ) : ( LB2D_shift_6 ) ;
assign n135 =  ( n30 ) ? ( LB2D_shift_6 ) : ( n134 ) ;
assign n136 =  ( n25 ) ? ( LB2D_shift_5 ) : ( n135 ) ;
assign n137 =  ( n18 ) ? ( LB2D_shift_6 ) : ( n136 ) ;
assign n138 =  ( n9 ) ? ( LB2D_shift_6 ) : ( n137 ) ;
assign n139 =  ( n4 ) ? ( LB2D_shift_6 ) : ( n138 ) ;
assign n140 =  ( n35 ) ? ( LB2D_shift_7 ) : ( LB2D_shift_7 ) ;
assign n141 =  ( n30 ) ? ( LB2D_shift_7 ) : ( n140 ) ;
assign n142 =  ( n25 ) ? ( LB2D_shift_6 ) : ( n141 ) ;
assign n143 =  ( n18 ) ? ( LB2D_shift_7 ) : ( n142 ) ;
assign n144 =  ( n9 ) ? ( LB2D_shift_7 ) : ( n143 ) ;
assign n145 =  ( n4 ) ? ( LB2D_shift_7 ) : ( n144 ) ;
assign n146 =  ( LB2D_shift_x ) + ( 9'd1 )  ;
assign n147 =  ( n35 ) ? ( LB2D_shift_x ) : ( LB2D_shift_x ) ;
assign n148 =  ( n30 ) ? ( LB2D_shift_x ) : ( n147 ) ;
assign n149 =  ( n25 ) ? ( n146 ) : ( n148 ) ;
assign n150 =  ( n18 ) ? ( LB2D_shift_x ) : ( n149 ) ;
assign n151 =  ( n9 ) ? ( LB2D_shift_x ) : ( n150 ) ;
assign n152 =  ( n4 ) ? ( LB2D_shift_x ) : ( n151 ) ;
assign n153 =  ( LB2D_shift_y ) < ( 10'd480 )  ;
assign n154 =  ( LB2D_shift_x ) < ( 9'd488 )  ;
assign n155 =  ( LB2D_shift_y ) + ( 10'd1 )  ;
assign n156 =  ( n154 ) ? ( LB2D_shift_y ) : ( n155 ) ;
assign n157 =  ( n153 ) ? ( n156 ) : ( 10'd480 ) ;
assign n158 =  ( n35 ) ? ( LB2D_shift_y ) : ( LB2D_shift_y ) ;
assign n159 =  ( n30 ) ? ( LB2D_shift_y ) : ( n158 ) ;
assign n160 =  ( n25 ) ? ( n157 ) : ( n159 ) ;
assign n161 =  ( n18 ) ? ( LB2D_shift_y ) : ( n160 ) ;
assign n162 =  ( n9 ) ? ( LB2D_shift_y ) : ( n161 ) ;
assign n163 =  ( n4 ) ? ( LB2D_shift_y ) : ( n162 ) ;
assign n164 =  ( stencil_stream_full ) == ( 1'd1 )  ;
assign n165 =  ( n164 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_0 ) ;
//assign n166 = gb_fun(n165) ;
gb_fun gb_fun_U (
        .a (n165),
        .b (n166)
        );
assign n167 =  ( n35 ) ? ( arg_0_TDATA ) : ( arg_0_TDATA ) ;
assign n168 =  ( n30 ) ? ( arg_0_TDATA ) : ( n167 ) ;
assign n169 =  ( n25 ) ? ( arg_0_TDATA ) : ( n168 ) ;
assign n170 =  ( n18 ) ? ( n166 ) : ( n169 ) ;
assign n171 =  ( n9 ) ? ( arg_0_TDATA ) : ( n170 ) ;
assign n172 =  ( n4 ) ? ( arg_0_TDATA ) : ( n171 ) ;
assign n173 =  ( gb_pp_it_8 ) == ( 1'd1 )  ;
assign n174 =  ( n173 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n175 =  ( n35 ) ? ( arg_0_TVALID ) : ( arg_0_TVALID ) ;
assign n176 =  ( n30 ) ? ( arg_0_TVALID ) : ( n175 ) ;
assign n177 =  ( n25 ) ? ( arg_0_TVALID ) : ( n176 ) ;
assign n178 =  ( n18 ) ? ( n174 ) : ( n177 ) ;
assign n179 =  ( n9 ) ? ( arg_0_TVALID ) : ( n178 ) ;
assign n180 =  ( n4 ) ? ( 1'd0 ) : ( n179 ) ;
assign n181 =  ( n35 ) ? ( 1'd1 ) : ( arg_1_TREADY ) ;
assign n182 =  ( n49 ) ? ( 1'd1 ) : ( n181 ) ;
assign n183 =  ( n30 ) ? ( arg_1_TREADY ) : ( n182 ) ;
assign n184 =  ( n25 ) ? ( arg_1_TREADY ) : ( n183 ) ;
assign n185 =  ( n18 ) ? ( arg_1_TREADY ) : ( n184 ) ;
assign n186 =  ( n9 ) ? ( 1'd0 ) : ( n185 ) ;
assign n187 =  ( n4 ) ? ( 1'd0 ) : ( n186 ) ;
assign n188 =  ( gb_p_cnt ) + ( 19'd1 )  ;
assign n189 =  ( n188 ) == ( 19'd307200 )  ;
assign n190 =  ( n189 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n191 =  ( n35 ) ? ( gb_exit_it_1 ) : ( gb_exit_it_1 ) ;
assign n192 =  ( n30 ) ? ( gb_exit_it_1 ) : ( n191 ) ;
assign n193 =  ( n25 ) ? ( gb_exit_it_1 ) : ( n192 ) ;
assign n194 =  ( n18 ) ? ( n190 ) : ( n193 ) ;
assign n195 =  ( n9 ) ? ( gb_exit_it_1 ) : ( n194 ) ;
assign n196 =  ( n4 ) ? ( gb_exit_it_1 ) : ( n195 ) ;
assign n197 =  ( n35 ) ? ( gb_exit_it_2 ) : ( gb_exit_it_2 ) ;
assign n198 =  ( n30 ) ? ( gb_exit_it_2 ) : ( n197 ) ;
assign n199 =  ( n25 ) ? ( gb_exit_it_2 ) : ( n198 ) ;
assign n200 =  ( n18 ) ? ( gb_exit_it_1 ) : ( n199 ) ;
assign n201 =  ( n9 ) ? ( gb_exit_it_2 ) : ( n200 ) ;
assign n202 =  ( n4 ) ? ( gb_exit_it_2 ) : ( n201 ) ;
assign n203 =  ( n35 ) ? ( gb_exit_it_3 ) : ( gb_exit_it_3 ) ;
assign n204 =  ( n30 ) ? ( gb_exit_it_3 ) : ( n203 ) ;
assign n205 =  ( n25 ) ? ( gb_exit_it_3 ) : ( n204 ) ;
assign n206 =  ( n18 ) ? ( gb_exit_it_2 ) : ( n205 ) ;
assign n207 =  ( n9 ) ? ( gb_exit_it_3 ) : ( n206 ) ;
assign n208 =  ( n4 ) ? ( gb_exit_it_3 ) : ( n207 ) ;
assign n209 =  ( n35 ) ? ( gb_exit_it_4 ) : ( gb_exit_it_4 ) ;
assign n210 =  ( n30 ) ? ( gb_exit_it_4 ) : ( n209 ) ;
assign n211 =  ( n25 ) ? ( gb_exit_it_4 ) : ( n210 ) ;
assign n212 =  ( n18 ) ? ( gb_exit_it_3 ) : ( n211 ) ;
assign n213 =  ( n9 ) ? ( gb_exit_it_4 ) : ( n212 ) ;
assign n214 =  ( n4 ) ? ( gb_exit_it_4 ) : ( n213 ) ;
assign n215 =  ( n35 ) ? ( gb_exit_it_5 ) : ( gb_exit_it_5 ) ;
assign n216 =  ( n30 ) ? ( gb_exit_it_5 ) : ( n215 ) ;
assign n217 =  ( n25 ) ? ( gb_exit_it_5 ) : ( n216 ) ;
assign n218 =  ( n18 ) ? ( gb_exit_it_4 ) : ( n217 ) ;
assign n219 =  ( n9 ) ? ( gb_exit_it_5 ) : ( n218 ) ;
assign n220 =  ( n4 ) ? ( gb_exit_it_5 ) : ( n219 ) ;
assign n221 =  ( n35 ) ? ( gb_exit_it_6 ) : ( gb_exit_it_6 ) ;
assign n222 =  ( n30 ) ? ( gb_exit_it_6 ) : ( n221 ) ;
assign n223 =  ( n25 ) ? ( gb_exit_it_6 ) : ( n222 ) ;
assign n224 =  ( n18 ) ? ( gb_exit_it_5 ) : ( n223 ) ;
assign n225 =  ( n9 ) ? ( gb_exit_it_6 ) : ( n224 ) ;
assign n226 =  ( n4 ) ? ( gb_exit_it_6 ) : ( n225 ) ;
assign n227 =  ( n35 ) ? ( gb_exit_it_7 ) : ( gb_exit_it_7 ) ;
assign n228 =  ( n30 ) ? ( gb_exit_it_7 ) : ( n227 ) ;
assign n229 =  ( n25 ) ? ( gb_exit_it_7 ) : ( n228 ) ;
assign n230 =  ( n18 ) ? ( gb_exit_it_6 ) : ( n229 ) ;
assign n231 =  ( n9 ) ? ( gb_exit_it_7 ) : ( n230 ) ;
assign n232 =  ( n4 ) ? ( gb_exit_it_7 ) : ( n231 ) ;
assign n233 =  ( n35 ) ? ( gb_exit_it_8 ) : ( gb_exit_it_8 ) ;
assign n234 =  ( n30 ) ? ( gb_exit_it_8 ) : ( n233 ) ;
assign n235 =  ( n25 ) ? ( gb_exit_it_8 ) : ( n234 ) ;
assign n236 =  ( n18 ) ? ( gb_exit_it_7 ) : ( n235 ) ;
assign n237 =  ( n9 ) ? ( gb_exit_it_8 ) : ( n236 ) ;
assign n238 =  ( n4 ) ? ( gb_exit_it_8 ) : ( n237 ) ;
assign n239 =  ( gb_p_cnt ) < ( 19'd307200 )  ;
assign n240 =  ( n239 ) ? ( n188 ) : ( 19'd307200 ) ;
assign n241 =  ( n35 ) ? ( gb_p_cnt ) : ( gb_p_cnt ) ;
assign n242 =  ( n30 ) ? ( gb_p_cnt ) : ( n241 ) ;
assign n243 =  ( n25 ) ? ( gb_p_cnt ) : ( n242 ) ;
assign n244 =  ( n18 ) ? ( n240 ) : ( n243 ) ;
assign n245 =  ( n9 ) ? ( gb_p_cnt ) : ( n244 ) ;
assign n246 =  ( n4 ) ? ( gb_p_cnt ) : ( n245 ) ;
assign n247 =  ( n35 ) ? ( gb_pp_it_1 ) : ( gb_pp_it_1 ) ;
assign n248 =  ( n30 ) ? ( gb_pp_it_1 ) : ( n247 ) ;
assign n249 =  ( n25 ) ? ( gb_pp_it_1 ) : ( n248 ) ;
assign n250 =  ( n18 ) ? ( 1'd1 ) : ( n249 ) ;
assign n251 =  ( n9 ) ? ( gb_pp_it_1 ) : ( n250 ) ;
assign n252 =  ( n4 ) ? ( gb_pp_it_1 ) : ( n251 ) ;
assign n253 =  ( n35 ) ? ( gb_pp_it_2 ) : ( gb_pp_it_2 ) ;
assign n254 =  ( n30 ) ? ( gb_pp_it_2 ) : ( n253 ) ;
assign n255 =  ( n25 ) ? ( gb_pp_it_2 ) : ( n254 ) ;
assign n256 =  ( n18 ) ? ( gb_pp_it_1 ) : ( n255 ) ;
assign n257 =  ( n9 ) ? ( gb_pp_it_2 ) : ( n256 ) ;
assign n258 =  ( n4 ) ? ( gb_pp_it_2 ) : ( n257 ) ;
assign n259 =  ( n35 ) ? ( gb_pp_it_3 ) : ( gb_pp_it_3 ) ;
assign n260 =  ( n30 ) ? ( gb_pp_it_3 ) : ( n259 ) ;
assign n261 =  ( n25 ) ? ( gb_pp_it_3 ) : ( n260 ) ;
assign n262 =  ( n18 ) ? ( gb_pp_it_2 ) : ( n261 ) ;
assign n263 =  ( n9 ) ? ( gb_pp_it_3 ) : ( n262 ) ;
assign n264 =  ( n4 ) ? ( gb_pp_it_3 ) : ( n263 ) ;
assign n265 =  ( n35 ) ? ( gb_pp_it_4 ) : ( gb_pp_it_4 ) ;
assign n266 =  ( n30 ) ? ( gb_pp_it_4 ) : ( n265 ) ;
assign n267 =  ( n25 ) ? ( gb_pp_it_4 ) : ( n266 ) ;
assign n268 =  ( n18 ) ? ( gb_pp_it_3 ) : ( n267 ) ;
assign n269 =  ( n9 ) ? ( gb_pp_it_4 ) : ( n268 ) ;
assign n270 =  ( n4 ) ? ( gb_pp_it_4 ) : ( n269 ) ;
assign n271 =  ( n35 ) ? ( gb_pp_it_5 ) : ( gb_pp_it_5 ) ;
assign n272 =  ( n30 ) ? ( gb_pp_it_5 ) : ( n271 ) ;
assign n273 =  ( n25 ) ? ( gb_pp_it_5 ) : ( n272 ) ;
assign n274 =  ( n18 ) ? ( gb_pp_it_4 ) : ( n273 ) ;
assign n275 =  ( n9 ) ? ( gb_pp_it_5 ) : ( n274 ) ;
assign n276 =  ( n4 ) ? ( gb_pp_it_5 ) : ( n275 ) ;
assign n277 =  ( n35 ) ? ( gb_pp_it_6 ) : ( gb_pp_it_6 ) ;
assign n278 =  ( n30 ) ? ( gb_pp_it_6 ) : ( n277 ) ;
assign n279 =  ( n25 ) ? ( gb_pp_it_6 ) : ( n278 ) ;
assign n280 =  ( n18 ) ? ( gb_pp_it_5 ) : ( n279 ) ;
assign n281 =  ( n9 ) ? ( gb_pp_it_6 ) : ( n280 ) ;
assign n282 =  ( n4 ) ? ( gb_pp_it_6 ) : ( n281 ) ;
assign n283 =  ( n35 ) ? ( gb_pp_it_7 ) : ( gb_pp_it_7 ) ;
assign n284 =  ( n30 ) ? ( gb_pp_it_7 ) : ( n283 ) ;
assign n285 =  ( n25 ) ? ( gb_pp_it_7 ) : ( n284 ) ;
assign n286 =  ( n18 ) ? ( gb_pp_it_6 ) : ( n285 ) ;
assign n287 =  ( n9 ) ? ( gb_pp_it_7 ) : ( n286 ) ;
assign n288 =  ( n4 ) ? ( gb_pp_it_7 ) : ( n287 ) ;
assign n289 =  ( n35 ) ? ( gb_pp_it_8 ) : ( gb_pp_it_8 ) ;
assign n290 =  ( n30 ) ? ( gb_pp_it_8 ) : ( n289 ) ;
assign n291 =  ( n25 ) ? ( gb_pp_it_8 ) : ( n290 ) ;
assign n292 =  ( n18 ) ? ( gb_pp_it_7 ) : ( n291 ) ;
assign n293 =  ( n9 ) ? ( gb_pp_it_8 ) : ( n292 ) ;
assign n294 =  ( n4 ) ? ( gb_pp_it_8 ) : ( n293 ) ;
assign n295 =  ( n35 ) ? ( gb_pp_it_9 ) : ( gb_pp_it_9 ) ;
assign n296 =  ( n30 ) ? ( gb_pp_it_9 ) : ( n295 ) ;
assign n297 =  ( n25 ) ? ( gb_pp_it_9 ) : ( n296 ) ;
assign n298 =  ( n18 ) ? ( gb_pp_it_8 ) : ( n297 ) ;
assign n299 =  ( n9 ) ? ( gb_pp_it_9 ) : ( n298 ) ;
assign n300 =  ( n4 ) ? ( gb_pp_it_9 ) : ( n299 ) ;
assign n301 =  ( n35 ) ? ( LB1D_buff ) : ( in_stream_buff_0 ) ;
assign n302 =  ( n30 ) ? ( in_stream_buff_0 ) : ( n301 ) ;
assign n303 =  ( n25 ) ? ( in_stream_buff_0 ) : ( n302 ) ;
assign n304 =  ( n18 ) ? ( in_stream_buff_0 ) : ( n303 ) ;
assign n305 =  ( n9 ) ? ( in_stream_buff_0 ) : ( n304 ) ;
assign n306 =  ( n4 ) ? ( in_stream_buff_0 ) : ( n305 ) ;
assign n307 =  ( n35 ) ? ( in_stream_buff_0 ) : ( in_stream_buff_1 ) ;
assign n308 =  ( n30 ) ? ( in_stream_buff_1 ) : ( n307 ) ;
assign n309 =  ( n25 ) ? ( in_stream_buff_1 ) : ( n308 ) ;
assign n310 =  ( n18 ) ? ( in_stream_buff_1 ) : ( n309 ) ;
assign n311 =  ( n9 ) ? ( in_stream_buff_1 ) : ( n310 ) ;
assign n312 =  ( n4 ) ? ( in_stream_buff_1 ) : ( n311 ) ;
assign n313 =  ( in_stream_full ) == ( 1'd1 )  ;
assign n314 =  ( n313 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n315 =  ( n35 ) ? ( 1'd0 ) : ( in_stream_empty ) ;
assign n316 =  ( n30 ) ? ( n314 ) : ( n315 ) ;
assign n317 =  ( n25 ) ? ( in_stream_empty ) : ( n316 ) ;
assign n318 =  ( n18 ) ? ( in_stream_empty ) : ( n317 ) ;
assign n319 =  ( n9 ) ? ( in_stream_empty ) : ( n318 ) ;
assign n320 =  ( n4 ) ? ( in_stream_empty ) : ( n319 ) ;
assign n321 =  ( in_stream_empty ) == ( 1'd1 )  ;
assign n322 =  ( n321 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n323 =  ( n35 ) ? ( n322 ) : ( in_stream_full ) ;
assign n324 =  ( n30 ) ? ( 1'd0 ) : ( n323 ) ;
assign n325 =  ( n25 ) ? ( in_stream_full ) : ( n324 ) ;
assign n326 =  ( n18 ) ? ( in_stream_full ) : ( n325 ) ;
assign n327 =  ( n9 ) ? ( in_stream_full ) : ( n326 ) ;
assign n328 =  ( n4 ) ? ( in_stream_full ) : ( n327 ) ;
assign n329 =  ( n313 ) ? ( in_stream_buff_1 ) : ( in_stream_buff_0 ) ;
assign n330 =  ( LB2D_proc_w ) == ( 64'd0 )  ;
assign n331 =  (  LB2D_proc_7 [ LB2D_proc_x ] )  ;
assign n332 =  ( LB2D_proc_w ) == ( 64'd1 )  ;
assign n333 =  (  LB2D_proc_0 [ LB2D_proc_x ] )  ;
assign n334 =  ( LB2D_proc_w ) == ( 64'd2 )  ;
assign n335 =  (  LB2D_proc_1 [ LB2D_proc_x ] )  ;
assign n336 =  ( LB2D_proc_w ) == ( 64'd3 )  ;
assign n337 =  (  LB2D_proc_2 [ LB2D_proc_x ] )  ;
assign n338 =  ( LB2D_proc_w ) == ( 64'd4 )  ;
assign n339 =  (  LB2D_proc_3 [ LB2D_proc_x ] )  ;
assign n340 =  ( LB2D_proc_w ) == ( 64'd5 )  ;
assign n341 =  (  LB2D_proc_4 [ LB2D_proc_x ] )  ;
assign n342 =  ( LB2D_proc_w ) == ( 64'd6 )  ;
assign n343 =  (  LB2D_proc_5 [ LB2D_proc_x ] )  ;
assign n344 =  (  LB2D_proc_6 [ LB2D_proc_x ] )  ;
assign n345 =  ( n342 ) ? ( n343 ) : ( n344 ) ;
assign n346 =  ( n340 ) ? ( n341 ) : ( n345 ) ;
assign n347 =  ( n338 ) ? ( n339 ) : ( n346 ) ;
assign n348 =  ( n336 ) ? ( n337 ) : ( n347 ) ;
assign n349 =  ( n334 ) ? ( n335 ) : ( n348 ) ;
assign n350 =  ( n332 ) ? ( n333 ) : ( n349 ) ;
assign n351 =  ( n330 ) ? ( n331 ) : ( n350 ) ;
assign n352 =  ( n342 ) ? ( n341 ) : ( n343 ) ;
assign n353 =  ( n340 ) ? ( n339 ) : ( n352 ) ;
assign n354 =  ( n338 ) ? ( n337 ) : ( n353 ) ;
assign n355 =  ( n336 ) ? ( n335 ) : ( n354 ) ;
assign n356 =  ( n334 ) ? ( n333 ) : ( n355 ) ;
assign n357 =  ( n332 ) ? ( n331 ) : ( n356 ) ;
assign n358 =  ( n330 ) ? ( n344 ) : ( n357 ) ;
assign n359 =  ( n342 ) ? ( n339 ) : ( n341 ) ;
assign n360 =  ( n340 ) ? ( n337 ) : ( n359 ) ;
assign n361 =  ( n338 ) ? ( n335 ) : ( n360 ) ;
assign n362 =  ( n336 ) ? ( n333 ) : ( n361 ) ;
assign n363 =  ( n334 ) ? ( n331 ) : ( n362 ) ;
assign n364 =  ( n332 ) ? ( n344 ) : ( n363 ) ;
assign n365 =  ( n330 ) ? ( n343 ) : ( n364 ) ;
assign n366 =  ( n342 ) ? ( n337 ) : ( n339 ) ;
assign n367 =  ( n340 ) ? ( n335 ) : ( n366 ) ;
assign n368 =  ( n338 ) ? ( n333 ) : ( n367 ) ;
assign n369 =  ( n336 ) ? ( n331 ) : ( n368 ) ;
assign n370 =  ( n334 ) ? ( n344 ) : ( n369 ) ;
assign n371 =  ( n332 ) ? ( n343 ) : ( n370 ) ;
assign n372 =  ( n330 ) ? ( n341 ) : ( n371 ) ;
assign n373 =  ( n342 ) ? ( n335 ) : ( n337 ) ;
assign n374 =  ( n340 ) ? ( n333 ) : ( n373 ) ;
assign n375 =  ( n338 ) ? ( n331 ) : ( n374 ) ;
assign n376 =  ( n336 ) ? ( n344 ) : ( n375 ) ;
assign n377 =  ( n334 ) ? ( n343 ) : ( n376 ) ;
assign n378 =  ( n332 ) ? ( n341 ) : ( n377 ) ;
assign n379 =  ( n330 ) ? ( n339 ) : ( n378 ) ;
assign n380 =  ( n342 ) ? ( n333 ) : ( n335 ) ;
assign n381 =  ( n340 ) ? ( n331 ) : ( n380 ) ;
assign n382 =  ( n338 ) ? ( n344 ) : ( n381 ) ;
assign n383 =  ( n336 ) ? ( n343 ) : ( n382 ) ;
assign n384 =  ( n334 ) ? ( n341 ) : ( n383 ) ;
assign n385 =  ( n332 ) ? ( n339 ) : ( n384 ) ;
assign n386 =  ( n330 ) ? ( n337 ) : ( n385 ) ;
assign n387 =  ( n342 ) ? ( n331 ) : ( n333 ) ;
assign n388 =  ( n340 ) ? ( n344 ) : ( n387 ) ;
assign n389 =  ( n338 ) ? ( n343 ) : ( n388 ) ;
assign n390 =  ( n336 ) ? ( n341 ) : ( n389 ) ;
assign n391 =  ( n334 ) ? ( n339 ) : ( n390 ) ;
assign n392 =  ( n332 ) ? ( n337 ) : ( n391 ) ;
assign n393 =  ( n330 ) ? ( n335 ) : ( n392 ) ;
assign n394 =  ( n342 ) ? ( n344 ) : ( n331 ) ;
assign n395 =  ( n340 ) ? ( n343 ) : ( n394 ) ;
assign n396 =  ( n338 ) ? ( n341 ) : ( n395 ) ;
assign n397 =  ( n336 ) ? ( n339 ) : ( n396 ) ;
assign n398 =  ( n334 ) ? ( n337 ) : ( n397 ) ;
assign n399 =  ( n332 ) ? ( n335 ) : ( n398 ) ;
assign n400 =  ( n330 ) ? ( n333 ) : ( n399 ) ;
assign n401 =  { ( n393 ) , ( n400 ) }  ;
assign n402 =  { ( n386 ) , ( n401 ) }  ;
assign n403 =  { ( n379 ) , ( n402 ) }  ;
assign n404 =  { ( n372 ) , ( n403 ) }  ;
assign n405 =  { ( n365 ) , ( n404 ) }  ;
assign n406 =  { ( n358 ) , ( n405 ) }  ;
assign n407 =  { ( n351 ) , ( n406 ) }  ;
assign n408 =  { ( n329 ) , ( n407 ) }  ;
assign n409 =  ( n28 ) ? ( slice_stream_buff_0 ) : ( n408 ) ;
assign n410 =  ( n35 ) ? ( slice_stream_buff_0 ) : ( slice_stream_buff_0 ) ;
assign n411 =  ( n30 ) ? ( n409 ) : ( n410 ) ;
assign n412 =  ( n25 ) ? ( slice_stream_buff_0 ) : ( n411 ) ;
assign n413 =  ( n18 ) ? ( slice_stream_buff_0 ) : ( n412 ) ;
assign n414 =  ( n9 ) ? ( slice_stream_buff_0 ) : ( n413 ) ;
assign n415 =  ( n4 ) ? ( slice_stream_buff_0 ) : ( n414 ) ;
assign n416 =  ( n28 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n417 =  ( n35 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_1 ) ;
assign n418 =  ( n30 ) ? ( n416 ) : ( n417 ) ;
assign n419 =  ( n25 ) ? ( slice_stream_buff_1 ) : ( n418 ) ;
assign n420 =  ( n18 ) ? ( slice_stream_buff_1 ) : ( n419 ) ;
assign n421 =  ( n9 ) ? ( slice_stream_buff_1 ) : ( n420 ) ;
assign n422 =  ( n4 ) ? ( slice_stream_buff_1 ) : ( n421 ) ;
assign n423 =  ( n96 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n424 =  ( n28 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n425 =  ( n35 ) ? ( slice_stream_empty ) : ( slice_stream_empty ) ;
assign n426 =  ( n30 ) ? ( n424 ) : ( n425 ) ;
assign n427 =  ( n25 ) ? ( n423 ) : ( n426 ) ;
assign n428 =  ( n18 ) ? ( slice_stream_empty ) : ( n427 ) ;
assign n429 =  ( n9 ) ? ( slice_stream_empty ) : ( n428 ) ;
assign n430 =  ( n4 ) ? ( slice_stream_empty ) : ( n429 ) ;
assign n431 =  ( slice_stream_empty ) == ( 1'd1 )  ;
assign n432 =  ( n431 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n433 =  ( n28 ) ? ( 1'd0 ) : ( n432 ) ;
assign n434 =  ( n35 ) ? ( slice_stream_full ) : ( slice_stream_full ) ;
assign n435 =  ( n30 ) ? ( n433 ) : ( n434 ) ;
assign n436 =  ( n25 ) ? ( 1'd0 ) : ( n435 ) ;
assign n437 =  ( n18 ) ? ( slice_stream_full ) : ( n436 ) ;
assign n438 =  ( n9 ) ? ( slice_stream_full ) : ( n437 ) ;
assign n439 =  ( n4 ) ? ( slice_stream_full ) : ( n438 ) ;
assign n440 =  ( LB2D_shift_x ) >= ( 9'd8 )  ;
assign n441 = n97[71:64] ;
assign n442 = LB2D_shift_0[71:64] ;
assign n443 = LB2D_shift_1[71:64] ;
assign n444 = LB2D_shift_2[71:64] ;
assign n445 = LB2D_shift_3[71:64] ;
assign n446 = LB2D_shift_4[71:64] ;
assign n447 = LB2D_shift_5[71:64] ;
assign n448 = LB2D_shift_6[71:64] ;
assign n449 = LB2D_shift_7[71:64] ;
assign n450 =  { ( n448 ) , ( n449 ) }  ;
assign n451 =  { ( n447 ) , ( n450 ) }  ;
assign n452 =  { ( n446 ) , ( n451 ) }  ;
assign n453 =  { ( n445 ) , ( n452 ) }  ;
assign n454 =  { ( n444 ) , ( n453 ) }  ;
assign n455 =  { ( n443 ) , ( n454 ) }  ;
assign n456 =  { ( n442 ) , ( n455 ) }  ;
assign n457 =  { ( n441 ) , ( n456 ) }  ;
assign n458 = n97[63:56] ;
assign n459 = LB2D_shift_0[63:56] ;
assign n460 = LB2D_shift_1[63:56] ;
assign n461 = LB2D_shift_2[63:56] ;
assign n462 = LB2D_shift_3[63:56] ;
assign n463 = LB2D_shift_4[63:56] ;
assign n464 = LB2D_shift_5[63:56] ;
assign n465 = LB2D_shift_6[63:56] ;
assign n466 = LB2D_shift_7[63:56] ;
assign n467 =  { ( n465 ) , ( n466 ) }  ;
assign n468 =  { ( n464 ) , ( n467 ) }  ;
assign n469 =  { ( n463 ) , ( n468 ) }  ;
assign n470 =  { ( n462 ) , ( n469 ) }  ;
assign n471 =  { ( n461 ) , ( n470 ) }  ;
assign n472 =  { ( n460 ) , ( n471 ) }  ;
assign n473 =  { ( n459 ) , ( n472 ) }  ;
assign n474 =  { ( n458 ) , ( n473 ) }  ;
assign n475 = n97[55:48] ;
assign n476 = LB2D_shift_0[55:48] ;
assign n477 = LB2D_shift_1[55:48] ;
assign n478 = LB2D_shift_2[55:48] ;
assign n479 = LB2D_shift_3[55:48] ;
assign n480 = LB2D_shift_4[55:48] ;
assign n481 = LB2D_shift_5[55:48] ;
assign n482 = LB2D_shift_6[55:48] ;
assign n483 = LB2D_shift_7[55:48] ;
assign n484 =  { ( n482 ) , ( n483 ) }  ;
assign n485 =  { ( n481 ) , ( n484 ) }  ;
assign n486 =  { ( n480 ) , ( n485 ) }  ;
assign n487 =  { ( n479 ) , ( n486 ) }  ;
assign n488 =  { ( n478 ) , ( n487 ) }  ;
assign n489 =  { ( n477 ) , ( n488 ) }  ;
assign n490 =  { ( n476 ) , ( n489 ) }  ;
assign n491 =  { ( n475 ) , ( n490 ) }  ;
assign n492 = n97[47:40] ;
assign n493 = LB2D_shift_0[47:40] ;
assign n494 = LB2D_shift_1[47:40] ;
assign n495 = LB2D_shift_2[47:40] ;
assign n496 = LB2D_shift_3[47:40] ;
assign n497 = LB2D_shift_4[47:40] ;
assign n498 = LB2D_shift_5[47:40] ;
assign n499 = LB2D_shift_6[47:40] ;
assign n500 = LB2D_shift_7[47:40] ;
assign n501 =  { ( n499 ) , ( n500 ) }  ;
assign n502 =  { ( n498 ) , ( n501 ) }  ;
assign n503 =  { ( n497 ) , ( n502 ) }  ;
assign n504 =  { ( n496 ) , ( n503 ) }  ;
assign n505 =  { ( n495 ) , ( n504 ) }  ;
assign n506 =  { ( n494 ) , ( n505 ) }  ;
assign n507 =  { ( n493 ) , ( n506 ) }  ;
assign n508 =  { ( n492 ) , ( n507 ) }  ;
assign n509 = n97[39:32] ;
assign n510 = LB2D_shift_0[39:32] ;
assign n511 = LB2D_shift_1[39:32] ;
assign n512 = LB2D_shift_2[39:32] ;
assign n513 = LB2D_shift_3[39:32] ;
assign n514 = LB2D_shift_4[39:32] ;
assign n515 = LB2D_shift_5[39:32] ;
assign n516 = LB2D_shift_6[39:32] ;
assign n517 = LB2D_shift_7[39:32] ;
assign n518 =  { ( n516 ) , ( n517 ) }  ;
assign n519 =  { ( n515 ) , ( n518 ) }  ;
assign n520 =  { ( n514 ) , ( n519 ) }  ;
assign n521 =  { ( n513 ) , ( n520 ) }  ;
assign n522 =  { ( n512 ) , ( n521 ) }  ;
assign n523 =  { ( n511 ) , ( n522 ) }  ;
assign n524 =  { ( n510 ) , ( n523 ) }  ;
assign n525 =  { ( n509 ) , ( n524 ) }  ;
assign n526 = n97[31:24] ;
assign n527 = LB2D_shift_0[31:24] ;
assign n528 = LB2D_shift_1[31:24] ;
assign n529 = LB2D_shift_2[31:24] ;
assign n530 = LB2D_shift_3[31:24] ;
assign n531 = LB2D_shift_4[31:24] ;
assign n532 = LB2D_shift_5[31:24] ;
assign n533 = LB2D_shift_6[31:24] ;
assign n534 = LB2D_shift_7[31:24] ;
assign n535 =  { ( n533 ) , ( n534 ) }  ;
assign n536 =  { ( n532 ) , ( n535 ) }  ;
assign n537 =  { ( n531 ) , ( n536 ) }  ;
assign n538 =  { ( n530 ) , ( n537 ) }  ;
assign n539 =  { ( n529 ) , ( n538 ) }  ;
assign n540 =  { ( n528 ) , ( n539 ) }  ;
assign n541 =  { ( n527 ) , ( n540 ) }  ;
assign n542 =  { ( n526 ) , ( n541 ) }  ;
assign n543 = n97[23:16] ;
assign n544 = LB2D_shift_0[23:16] ;
assign n545 = LB2D_shift_1[23:16] ;
assign n546 = LB2D_shift_2[23:16] ;
assign n547 = LB2D_shift_3[23:16] ;
assign n548 = LB2D_shift_4[23:16] ;
assign n549 = LB2D_shift_5[23:16] ;
assign n550 = LB2D_shift_6[23:16] ;
assign n551 = LB2D_shift_7[23:16] ;
assign n552 =  { ( n550 ) , ( n551 ) }  ;
assign n553 =  { ( n549 ) , ( n552 ) }  ;
assign n554 =  { ( n548 ) , ( n553 ) }  ;
assign n555 =  { ( n547 ) , ( n554 ) }  ;
assign n556 =  { ( n546 ) , ( n555 ) }  ;
assign n557 =  { ( n545 ) , ( n556 ) }  ;
assign n558 =  { ( n544 ) , ( n557 ) }  ;
assign n559 =  { ( n543 ) , ( n558 ) }  ;
assign n560 = n97[15:8] ;
assign n561 = LB2D_shift_0[15:8] ;
assign n562 = LB2D_shift_1[15:8] ;
assign n563 = LB2D_shift_2[15:8] ;
assign n564 = LB2D_shift_3[15:8] ;
assign n565 = LB2D_shift_4[15:8] ;
assign n566 = LB2D_shift_5[15:8] ;
assign n567 = LB2D_shift_6[15:8] ;
assign n568 = LB2D_shift_7[15:8] ;
assign n569 =  { ( n567 ) , ( n568 ) }  ;
assign n570 =  { ( n566 ) , ( n569 ) }  ;
assign n571 =  { ( n565 ) , ( n570 ) }  ;
assign n572 =  { ( n564 ) , ( n571 ) }  ;
assign n573 =  { ( n563 ) , ( n572 ) }  ;
assign n574 =  { ( n562 ) , ( n573 ) }  ;
assign n575 =  { ( n561 ) , ( n574 ) }  ;
assign n576 =  { ( n560 ) , ( n575 ) }  ;
assign n577 = n97[7:0] ;
assign n578 = LB2D_shift_0[7:0] ;
assign n579 = LB2D_shift_1[7:0] ;
assign n580 = LB2D_shift_2[7:0] ;
assign n581 = LB2D_shift_3[7:0] ;
assign n582 = LB2D_shift_4[7:0] ;
assign n583 = LB2D_shift_5[7:0] ;
assign n584 = LB2D_shift_6[7:0] ;
assign n585 = LB2D_shift_7[7:0] ;
assign n586 =  { ( n584 ) , ( n585 ) }  ;
assign n587 =  { ( n583 ) , ( n586 ) }  ;
assign n588 =  { ( n582 ) , ( n587 ) }  ;
assign n589 =  { ( n581 ) , ( n588 ) }  ;
assign n590 =  { ( n580 ) , ( n589 ) }  ;
assign n591 =  { ( n579 ) , ( n590 ) }  ;
assign n592 =  { ( n578 ) , ( n591 ) }  ;
assign n593 =  { ( n577 ) , ( n592 ) }  ;
assign n594 =  { ( n576 ) , ( n593 ) }  ;
assign n595 =  { ( n559 ) , ( n594 ) }  ;
assign n596 =  { ( n542 ) , ( n595 ) }  ;
assign n597 =  { ( n525 ) , ( n596 ) }  ;
assign n598 =  { ( n508 ) , ( n597 ) }  ;
assign n599 =  { ( n491 ) , ( n598 ) }  ;
assign n600 =  { ( n474 ) , ( n599 ) }  ;
assign n601 =  { ( n457 ) , ( n600 ) }  ;
assign n602 =  ( n440 ) ? ( n601 ) : ( stencil_stream_buff_0 ) ;
assign n603 =  ( n35 ) ? ( stencil_stream_buff_0 ) : ( stencil_stream_buff_0 ) ;
assign n604 =  ( n30 ) ? ( stencil_stream_buff_0 ) : ( n603 ) ;
assign n605 =  ( n25 ) ? ( n602 ) : ( n604 ) ;
assign n606 =  ( n18 ) ? ( stencil_stream_buff_0 ) : ( n605 ) ;
assign n607 =  ( n9 ) ? ( stencil_stream_buff_0 ) : ( n606 ) ;
assign n608 =  ( n4 ) ? ( stencil_stream_buff_0 ) : ( n607 ) ;
assign n609 =  ( n35 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_1 ) ;
assign n610 =  ( n30 ) ? ( stencil_stream_buff_1 ) : ( n609 ) ;
assign n611 =  ( n25 ) ? ( stencil_stream_buff_0 ) : ( n610 ) ;
assign n612 =  ( n18 ) ? ( stencil_stream_buff_1 ) : ( n611 ) ;
assign n613 =  ( n9 ) ? ( stencil_stream_buff_1 ) : ( n612 ) ;
assign n614 =  ( n4 ) ? ( stencil_stream_buff_1 ) : ( n613 ) ;
assign n615 =  ( n164 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n616 =  ( n23 ) ? ( stencil_stream_empty ) : ( 1'd0 ) ;
assign n617 =  ( n35 ) ? ( stencil_stream_empty ) : ( stencil_stream_empty ) ;
assign n618 =  ( n30 ) ? ( stencil_stream_empty ) : ( n617 ) ;
assign n619 =  ( n25 ) ? ( n616 ) : ( n618 ) ;
assign n620 =  ( n18 ) ? ( n615 ) : ( n619 ) ;
assign n621 =  ( n9 ) ? ( stencil_stream_empty ) : ( n620 ) ;
assign n622 =  ( n4 ) ? ( stencil_stream_empty ) : ( n621 ) ;
assign n623 =  ( n14 ) ? ( 1'd0 ) : ( 1'd0 ) ;
assign n624 =  ( stencil_stream_empty ) == ( 1'd1 )  ;
assign n625 =  ( n624 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n626 =  ( n23 ) ? ( stencil_stream_full ) : ( n625 ) ;
assign n627 =  ( n35 ) ? ( stencil_stream_full ) : ( stencil_stream_full ) ;
assign n628 =  ( n30 ) ? ( stencil_stream_full ) : ( n627 ) ;
assign n629 =  ( n25 ) ? ( n626 ) : ( n628 ) ;
assign n630 =  ( n18 ) ? ( n623 ) : ( n629 ) ;
assign n631 =  ( n9 ) ? ( stencil_stream_full ) : ( n630 ) ;
assign n632 =  ( n4 ) ? ( stencil_stream_full ) : ( n631 ) ;
assign n633 = ~ ( n4 ) ;
assign n634 = ~ ( n9 ) ;
assign n635 =  ( n633 ) & ( n634 )  ;
assign n636 = ~ ( n18 ) ;
assign n637 =  ( n635 ) & ( n636 )  ;
assign n638 = ~ ( n25 ) ;
assign n639 =  ( n637 ) & ( n638 )  ;
assign n640 = ~ ( n30 ) ;
assign n641 =  ( n639 ) & ( n640 )  ;
assign n642 = ~ ( n35 ) ;
assign n643 =  ( n641 ) & ( n642 )  ;
assign n644 =  ( n641 ) & ( n35 )  ;
assign n645 =  ( n639 ) & ( n30 )  ;
assign n646 = ~ ( n330 ) ;
assign n647 =  ( n645 ) & ( n646 )  ;
assign n648 =  ( n645 ) & ( n330 )  ;
assign n649 =  ( n637 ) & ( n25 )  ;
assign n650 =  ( n635 ) & ( n18 )  ;
assign n651 =  ( n633 ) & ( n9 )  ;
assign LB2D_proc_0_addr0 = n648 ? (LB2D_proc_x) : (0);
assign LB2D_proc_0_data0 = n648 ? (n329) : (LB2D_proc_0[0]);
assign n652 = ~ ( n332 ) ;
assign n653 =  ( n645 ) & ( n652 )  ;
assign n654 =  ( n645 ) & ( n332 )  ;
assign LB2D_proc_1_addr0 = n654 ? (LB2D_proc_x) : (0);
assign LB2D_proc_1_data0 = n654 ? (n329) : (LB2D_proc_1[0]);
assign n655 = ~ ( n334 ) ;
assign n656 =  ( n645 ) & ( n655 )  ;
assign n657 =  ( n645 ) & ( n334 )  ;
assign LB2D_proc_2_addr0 = n657 ? (LB2D_proc_x) : (0);
assign LB2D_proc_2_data0 = n657 ? (n329) : (LB2D_proc_2[0]);
assign n658 = ~ ( n336 ) ;
assign n659 =  ( n645 ) & ( n658 )  ;
assign n660 =  ( n645 ) & ( n336 )  ;
assign LB2D_proc_3_addr0 = n660 ? (LB2D_proc_x) : (0);
assign LB2D_proc_3_data0 = n660 ? (n329) : (LB2D_proc_3[0]);
assign n661 = ~ ( n338 ) ;
assign n662 =  ( n645 ) & ( n661 )  ;
assign n663 =  ( n645 ) & ( n338 )  ;
assign LB2D_proc_4_addr0 = n663 ? (LB2D_proc_x) : (0);
assign LB2D_proc_4_data0 = n663 ? (n329) : (LB2D_proc_4[0]);
assign n664 = ~ ( n340 ) ;
assign n665 =  ( n645 ) & ( n664 )  ;
assign n666 =  ( n645 ) & ( n340 )  ;
assign LB2D_proc_5_addr0 = n666 ? (LB2D_proc_x) : (0);
assign LB2D_proc_5_data0 = n666 ? (n329) : (LB2D_proc_5[0]);
assign n667 = ~ ( n342 ) ;
assign n668 =  ( n645 ) & ( n667 )  ;
assign n669 =  ( n645 ) & ( n342 )  ;
assign LB2D_proc_6_addr0 = n669 ? (LB2D_proc_x) : (0);
assign LB2D_proc_6_data0 = n669 ? (n329) : (LB2D_proc_6[0]);
assign n670 = ~ ( n68 ) ;
assign n671 =  ( n645 ) & ( n670 )  ;
assign n672 =  ( n645 ) & ( n68 )  ;
assign LB2D_proc_7_addr0 = n672 ? (LB2D_proc_x) : (0);
assign LB2D_proc_7_data0 = n672 ? (n329) : (LB2D_proc_7[0]);
/*
function [7:0] gb_fun ;
input [647:0] arg0;
    begin
//TODO: Add the specific function HERE.    end
endfunction
*/

always @(posedge clk) begin
   if(rst) begin
       LB1D_buff <= LB1D_buff;
       LB1D_in <= LB1D_in;
       LB1D_it_1 <= LB1D_it_1;
       LB1D_p_cnt <= LB1D_p_cnt;
       LB1D_uIn <= LB1D_uIn;
       LB2D_proc_w <= LB2D_proc_w;
       LB2D_proc_x <= LB2D_proc_x;
       LB2D_proc_y <= LB2D_proc_y;
       LB2D_shift_0 <= LB2D_shift_0;
       LB2D_shift_1 <= LB2D_shift_1;
       LB2D_shift_2 <= LB2D_shift_2;
       LB2D_shift_3 <= LB2D_shift_3;
       LB2D_shift_4 <= LB2D_shift_4;
       LB2D_shift_5 <= LB2D_shift_5;
       LB2D_shift_6 <= LB2D_shift_6;
       LB2D_shift_7 <= LB2D_shift_7;
       LB2D_shift_x <= LB2D_shift_x;
       LB2D_shift_y <= LB2D_shift_y;
       arg_0_TDATA <= arg_0_TDATA;
       arg_0_TVALID <= arg_0_TVALID;
       arg_1_TREADY <= arg_1_TREADY;
       gb_exit_it_1 <= gb_exit_it_1;
       gb_exit_it_2 <= gb_exit_it_2;
       gb_exit_it_3 <= gb_exit_it_3;
       gb_exit_it_4 <= gb_exit_it_4;
       gb_exit_it_5 <= gb_exit_it_5;
       gb_exit_it_6 <= gb_exit_it_6;
       gb_exit_it_7 <= gb_exit_it_7;
       gb_exit_it_8 <= gb_exit_it_8;
       gb_p_cnt <= gb_p_cnt;
       gb_pp_it_1 <= gb_pp_it_1;
       gb_pp_it_2 <= gb_pp_it_2;
       gb_pp_it_3 <= gb_pp_it_3;
       gb_pp_it_4 <= gb_pp_it_4;
       gb_pp_it_5 <= gb_pp_it_5;
       gb_pp_it_6 <= gb_pp_it_6;
       gb_pp_it_7 <= gb_pp_it_7;
       gb_pp_it_8 <= gb_pp_it_8;
       gb_pp_it_9 <= gb_pp_it_9;
       in_stream_buff_0 <= in_stream_buff_0;
       in_stream_buff_1 <= in_stream_buff_1;
       in_stream_empty <= in_stream_empty;
       in_stream_full <= in_stream_full;
       slice_stream_buff_0 <= slice_stream_buff_0;
       slice_stream_buff_1 <= slice_stream_buff_1;
       slice_stream_empty <= slice_stream_empty;
       slice_stream_full <= slice_stream_full;
       stencil_stream_buff_0 <= stencil_stream_buff_0;
       stencil_stream_buff_1 <= stencil_stream_buff_1;
       stencil_stream_empty <= stencil_stream_empty;
       stencil_stream_full <= stencil_stream_full;
   end
   else if(step) begin
       LB1D_buff <= n41;
       LB1D_in <= n47;
       LB1D_it_1 <= n50;
       LB1D_p_cnt <= n61;
       LB1D_uIn <= n66;
       LB2D_proc_w <= n77;
       LB2D_proc_x <= n85;
       LB2D_proc_y <= n95;
       LB2D_shift_0 <= n103;
       LB2D_shift_1 <= n109;
       LB2D_shift_2 <= n115;
       LB2D_shift_3 <= n121;
       LB2D_shift_4 <= n127;
       LB2D_shift_5 <= n133;
       LB2D_shift_6 <= n139;
       LB2D_shift_7 <= n145;
       LB2D_shift_x <= n152;
       LB2D_shift_y <= n163;
       arg_0_TDATA <= n172;
       arg_0_TVALID <= n180;
       arg_1_TREADY <= n187;
       gb_exit_it_1 <= n196;
       gb_exit_it_2 <= n202;
       gb_exit_it_3 <= n208;
       gb_exit_it_4 <= n214;
       gb_exit_it_5 <= n220;
       gb_exit_it_6 <= n226;
       gb_exit_it_7 <= n232;
       gb_exit_it_8 <= n238;
       gb_p_cnt <= n246;
       gb_pp_it_1 <= n252;
       gb_pp_it_2 <= n258;
       gb_pp_it_3 <= n264;
       gb_pp_it_4 <= n270;
       gb_pp_it_5 <= n276;
       gb_pp_it_6 <= n282;
       gb_pp_it_7 <= n288;
       gb_pp_it_8 <= n294;
       gb_pp_it_9 <= n300;
       in_stream_buff_0 <= n306;
       in_stream_buff_1 <= n312;
       in_stream_empty <= n320;
       in_stream_full <= n328;
       slice_stream_buff_0 <= n415;
       slice_stream_buff_1 <= n422;
       slice_stream_empty <= n430;
       slice_stream_full <= n439;
       stencil_stream_buff_0 <= n608;
       stencil_stream_buff_1 <= n614;
       stencil_stream_empty <= n622;
       stencil_stream_full <= n632;
       LB2D_proc_0 [ LB2D_proc_0_addr0 ] <= LB2D_proc_0_data0;
       LB2D_proc_1 [ LB2D_proc_1_addr0 ] <= LB2D_proc_1_data0;
       LB2D_proc_2 [ LB2D_proc_2_addr0 ] <= LB2D_proc_2_data0;
       LB2D_proc_3 [ LB2D_proc_3_addr0 ] <= LB2D_proc_3_data0;
       LB2D_proc_4 [ LB2D_proc_4_addr0 ] <= LB2D_proc_4_data0;
       LB2D_proc_5 [ LB2D_proc_5_addr0 ] <= LB2D_proc_5_data0;
       LB2D_proc_6 [ LB2D_proc_6_addr0 ] <= LB2D_proc_6_data0;
       LB2D_proc_7 [ LB2D_proc_7_addr0 ] <= LB2D_proc_7_data0;
   end
end
endmodule
