/* PREHEADER */
module fun_gb_fun (
    input [647:0] arg1,
    output [7:0] result
);
//TODO: Add the specific function HERE.
endmodule

/* END OF PREHEADER */
module SPEC_A(
arg_0_TREADY,
arg_1_TDATA,
arg_1_TVALID,
RAM_w,
RAM_x,
RAM_y,
arg_0_TDATA,
arg_0_TVALID,
arg_1_TREADY,
cur_pix,
gbit,
pre_pix,
proc_in,
st_ready,
stencil_0,
stencil_1,
stencil_2,
stencil_3,
stencil_4,
stencil_5,
stencil_6,
stencil_7,
stencil_8,
clk,rst,
step
);
input            arg_0_TREADY;
input      [7:0] arg_1_TDATA;
input            arg_1_TVALID;
input clk;
input rst;
input step;
output      [2:0] RAM_w;
output      [8:0] RAM_x;
output      [9:0] RAM_y;
output      [7:0] arg_0_TDATA;
output            arg_0_TVALID;
output            arg_1_TREADY;
output      [7:0] cur_pix;
output      [3:0] gbit;
output      [7:0] pre_pix;
output    [647:0] proc_in;
output            st_ready;
output     [71:0] stencil_0;
output     [71:0] stencil_1;
output     [71:0] stencil_2;
output     [71:0] stencil_3;
output     [71:0] stencil_4;
output     [71:0] stencil_5;
output     [71:0] stencil_6;
output     [71:0] stencil_7;
output     [71:0] stencil_8;
reg      [2:0] RAM_w;
reg      [8:0] RAM_x;
reg      [9:0] RAM_y;
reg      [7:0] arg_0_TDATA;
reg            arg_0_TVALID;
reg            arg_1_TREADY;
reg      [7:0] cur_pix;
reg      [3:0] gbit;
reg      [7:0] pre_pix;
reg    [647:0] proc_in;
reg            st_ready;
reg     [71:0] stencil_0;
reg     [71:0] stencil_1;
reg     [71:0] stencil_2;
reg     [71:0] stencil_3;
reg     [71:0] stencil_4;
reg     [71:0] stencil_5;
reg     [71:0] stencil_6;
reg     [71:0] stencil_7;
reg     [71:0] stencil_8;
wire            arg_0_TREADY;
wire      [7:0] arg_1_TDATA;
wire            arg_1_TVALID;
wire            n0;
wire            n1;
wire            n2;
wire            n3;
wire            n4;
wire            n5;
wire            n6;
wire            n7;
wire            n8;
wire            n9;
wire            n10;
wire            n11;
wire            n12;
wire            n13;
wire      [2:0] n14;
wire      [2:0] n15;
wire      [2:0] n16;
wire            n17;
wire            n18;
wire            n19;
wire            n20;
wire            n21;
wire            n22;
wire      [2:0] n23;
wire      [2:0] n24;
wire      [2:0] n25;
wire      [2:0] n26;
wire            n27;
wire            n28;
wire            n29;
wire      [8:0] n30;
wire      [8:0] n31;
wire      [8:0] n32;
wire      [8:0] n33;
wire      [8:0] n34;
wire      [8:0] n35;
wire      [8:0] n36;
wire            n37;
wire      [9:0] n38;
wire      [9:0] n39;
wire      [9:0] n40;
wire      [9:0] n41;
wire      [9:0] n42;
wire      [9:0] n43;
wire      [9:0] n44;
wire            n45;
wire            n46;
wire            n47;
wire            n48;
wire            n49;
wire            n50;
wire            n51;
wire            n52;
wire      [7:0] n53;
wire      [7:0] n54;
wire      [7:0] n55;
wire      [7:0] n56;
wire      [7:0] n57;
wire      [7:0] n58;
wire      [7:0] n59;
wire      [7:0] n60;
wire      [7:0] n61;
wire     [15:0] n62;
wire     [23:0] n63;
wire     [31:0] n64;
wire     [39:0] n65;
wire     [47:0] n66;
wire     [55:0] n67;
wire     [63:0] n68;
wire     [71:0] n69;
wire      [7:0] n70;
wire      [7:0] n71;
wire      [7:0] n72;
wire      [7:0] n73;
wire      [7:0] n74;
wire      [7:0] n75;
wire      [7:0] n76;
wire      [7:0] n77;
wire      [7:0] n78;
wire     [15:0] n79;
wire     [23:0] n80;
wire     [31:0] n81;
wire     [39:0] n82;
wire     [47:0] n83;
wire     [55:0] n84;
wire     [63:0] n85;
wire     [71:0] n86;
wire      [7:0] n87;
wire      [7:0] n88;
wire      [7:0] n89;
wire      [7:0] n90;
wire      [7:0] n91;
wire      [7:0] n92;
wire      [7:0] n93;
wire      [7:0] n94;
wire      [7:0] n95;
wire     [15:0] n96;
wire     [23:0] n97;
wire     [31:0] n98;
wire     [39:0] n99;
wire     [47:0] n100;
wire     [55:0] n101;
wire     [63:0] n102;
wire     [71:0] n103;
wire      [7:0] n104;
wire      [7:0] n105;
wire      [7:0] n106;
wire      [7:0] n107;
wire      [7:0] n108;
wire      [7:0] n109;
wire      [7:0] n110;
wire      [7:0] n111;
wire      [7:0] n112;
wire     [15:0] n113;
wire     [23:0] n114;
wire     [31:0] n115;
wire     [39:0] n116;
wire     [47:0] n117;
wire     [55:0] n118;
wire     [63:0] n119;
wire     [71:0] n120;
wire      [7:0] n121;
wire      [7:0] n122;
wire      [7:0] n123;
wire      [7:0] n124;
wire      [7:0] n125;
wire      [7:0] n126;
wire      [7:0] n127;
wire      [7:0] n128;
wire      [7:0] n129;
wire     [15:0] n130;
wire     [23:0] n131;
wire     [31:0] n132;
wire     [39:0] n133;
wire     [47:0] n134;
wire     [55:0] n135;
wire     [63:0] n136;
wire     [71:0] n137;
wire      [7:0] n138;
wire      [7:0] n139;
wire      [7:0] n140;
wire      [7:0] n141;
wire      [7:0] n142;
wire      [7:0] n143;
wire      [7:0] n144;
wire      [7:0] n145;
wire      [7:0] n146;
wire     [15:0] n147;
wire     [23:0] n148;
wire     [31:0] n149;
wire     [39:0] n150;
wire     [47:0] n151;
wire     [55:0] n152;
wire     [63:0] n153;
wire     [71:0] n154;
wire      [7:0] n155;
wire      [7:0] n156;
wire      [7:0] n157;
wire      [7:0] n158;
wire      [7:0] n159;
wire      [7:0] n160;
wire      [7:0] n161;
wire      [7:0] n162;
wire      [7:0] n163;
wire     [15:0] n164;
wire     [23:0] n165;
wire     [31:0] n166;
wire     [39:0] n167;
wire     [47:0] n168;
wire     [55:0] n169;
wire     [63:0] n170;
wire     [71:0] n171;
wire      [7:0] n172;
wire      [7:0] n173;
wire      [7:0] n174;
wire      [7:0] n175;
wire      [7:0] n176;
wire      [7:0] n177;
wire      [7:0] n178;
wire      [7:0] n179;
wire      [7:0] n180;
wire     [15:0] n181;
wire     [23:0] n182;
wire     [31:0] n183;
wire     [39:0] n184;
wire     [47:0] n185;
wire     [55:0] n186;
wire     [63:0] n187;
wire     [71:0] n188;
wire      [7:0] n189;
wire      [7:0] n190;
wire      [7:0] n191;
wire      [7:0] n192;
wire      [7:0] n193;
wire      [7:0] n194;
wire      [7:0] n195;
wire      [7:0] n196;
wire      [7:0] n197;
wire     [15:0] n198;
wire     [23:0] n199;
wire     [31:0] n200;
wire     [39:0] n201;
wire     [47:0] n202;
wire     [55:0] n203;
wire     [63:0] n204;
wire     [71:0] n205;
wire    [143:0] n206;
wire    [215:0] n207;
wire    [287:0] n208;
wire    [359:0] n209;
wire    [431:0] n210;
wire    [503:0] n211;
wire    [575:0] n212;
wire    [647:0] n213;
wire    [647:0] n214;
wire    [647:0] n215;
wire      [7:0] n216;
wire      [7:0] n218;
wire      [7:0] n219;
wire      [7:0] n220;
wire      [7:0] n221;
wire      [7:0] n222;
wire      [7:0] n223;
wire            n224;
wire            n225;
wire            n226;
wire            n227;
wire            n228;
wire            n229;
wire            n230;
wire            n231;
wire            n232;
wire            n233;
wire            n234;
wire      [8:0] n235;
wire            n236;
wire      [9:0] n237;
wire            n238;
wire            n239;
wire            n240;
wire            n241;
wire            n242;
wire            n243;
wire            n244;
wire            n245;
wire            n246;
wire            n247;
wire      [7:0] n248;
wire      [7:0] n249;
wire      [7:0] n250;
wire      [7:0] n251;
wire            n252;
wire      [3:0] n253;
wire      [3:0] n254;
wire      [3:0] n255;
wire      [7:0] n256;
wire      [7:0] n257;
wire    [647:0] n258;
wire    [647:0] n259;
wire            n260;
wire            n261;
wire     [71:0] n262;
wire     [71:0] n263;
wire     [71:0] n264;
wire     [71:0] n265;
wire     [71:0] n266;
wire     [71:0] n267;
wire     [71:0] n268;
wire     [71:0] n269;
wire     [71:0] n270;
wire     [71:0] n271;
wire     [71:0] n272;
wire     [71:0] n273;
wire     [71:0] n274;
wire     [71:0] n275;
wire     [71:0] n276;
wire     [71:0] n277;
wire     [71:0] n278;
wire     [71:0] n279;
wire     [71:0] n280;
wire     [71:0] n281;
wire     [71:0] n282;
wire     [71:0] n283;
wire     [71:0] n284;
wire     [71:0] n285;
wire     [71:0] n286;
wire     [71:0] n287;
wire     [71:0] n288;
wire     [71:0] n289;
wire     [71:0] n290;
wire     [71:0] n291;
wire     [71:0] n292;
wire     [71:0] n293;
wire     [71:0] n294;
wire     [71:0] n295;
wire     [71:0] n296;
wire     [71:0] n297;
wire     [71:0] n298;
wire     [71:0] n299;
wire     [71:0] n300;
wire     [71:0] n301;
wire            n302;
wire      [8:0] n303;
wire      [7:0] n304;
wire            n305;
wire      [7:0] n306;
wire            n307;
wire      [7:0] n308;
wire            n309;
wire      [7:0] n310;
wire            n311;
wire      [7:0] n312;
wire            n313;
wire      [7:0] n314;
wire            n315;
wire      [7:0] n316;
wire      [7:0] n317;
wire      [7:0] n318;
wire      [7:0] n319;
wire      [7:0] n320;
wire      [7:0] n321;
wire      [7:0] n322;
wire      [7:0] n323;
wire      [7:0] n324;
wire      [7:0] n325;
wire      [7:0] n326;
wire      [7:0] n327;
wire      [7:0] n328;
wire      [7:0] n329;
wire      [7:0] n330;
wire      [7:0] n331;
wire      [7:0] n332;
wire      [7:0] n333;
wire      [7:0] n334;
wire      [7:0] n335;
wire      [7:0] n336;
wire      [7:0] n337;
wire      [7:0] n338;
wire      [7:0] n339;
wire      [7:0] n340;
wire      [7:0] n341;
wire      [7:0] n342;
wire      [7:0] n343;
wire      [7:0] n344;
wire      [7:0] n345;
wire      [7:0] n346;
wire      [7:0] n347;
wire      [7:0] n348;
wire      [7:0] n349;
wire      [7:0] n350;
wire      [7:0] n351;
wire      [7:0] n352;
wire      [7:0] n353;
wire      [7:0] n354;
wire      [7:0] n355;
wire      [7:0] n356;
wire      [7:0] n357;
wire      [7:0] n358;
wire      [7:0] n359;
wire      [7:0] n360;
wire      [7:0] n361;
wire      [7:0] n362;
wire      [7:0] n363;
wire      [7:0] n364;
wire      [7:0] n365;
wire      [7:0] n366;
wire      [7:0] n367;
wire      [7:0] n368;
wire      [7:0] n369;
wire      [7:0] n370;
wire      [7:0] n371;
wire      [7:0] n372;
wire      [7:0] n373;
wire     [15:0] n374;
wire     [23:0] n375;
wire     [31:0] n376;
wire     [39:0] n377;
wire     [47:0] n378;
wire     [55:0] n379;
wire     [63:0] n380;
wire     [71:0] n381;
wire     [71:0] n382;
wire     [71:0] n383;
wire     [71:0] n384;
wire     [71:0] n385;
wire     [71:0] n386;
wire      [8:0] RAM_0_addr0;
wire      [7:0] RAM_0_data0;
wire            RAM_0_wen0;
wire            n387;
wire            n388;
wire            n389;
wire            n390;
wire            n391;
wire            n392;
wire            n393;
wire            n394;
wire            n395;
wire            n396;
wire            n397;
wire            n398;
wire            n399;
wire            n400;
wire            n401;
wire            n402;
wire            n403;
wire            n404;
wire      [8:0] RAM_1_addr0;
wire      [7:0] RAM_1_data0;
wire            RAM_1_wen0;
wire            n405;
wire            n406;
wire            n407;
wire      [8:0] RAM_2_addr0;
wire      [7:0] RAM_2_data0;
wire            RAM_2_wen0;
wire            n408;
wire            n409;
wire            n410;
wire      [8:0] RAM_3_addr0;
wire      [7:0] RAM_3_data0;
wire            RAM_3_wen0;
wire            n411;
wire            n412;
wire            n413;
wire      [8:0] RAM_4_addr0;
wire      [7:0] RAM_4_data0;
wire            RAM_4_wen0;
wire            n414;
wire            n415;
wire            n416;
wire      [8:0] RAM_5_addr0;
wire      [7:0] RAM_5_data0;
wire            RAM_5_wen0;
wire            n417;
wire            n418;
wire            n419;
wire      [8:0] RAM_6_addr0;
wire      [7:0] RAM_6_data0;
wire            RAM_6_wen0;
wire            n420;
wire            n421;
wire            n422;
wire      [8:0] RAM_7_addr0;
wire      [7:0] RAM_7_data0;
wire            RAM_7_wen0;
wire            n423;
wire            n424;
wire            n425;
reg      [7:0] RAM_0[511:0];
reg      [7:0] RAM_1[511:0];
reg      [7:0] RAM_2[511:0];
reg      [7:0] RAM_3[511:0];
reg      [7:0] RAM_4[511:0];
reg      [7:0] RAM_5[511:0];
reg      [7:0] RAM_6[511:0];
reg      [7:0] RAM_7[511:0];
wire clk;
wire rst;
wire step;
assign n0 =  ( arg_1_TVALID ) == ( 1'd0 )  ;
assign n1 =  ( arg_0_TVALID ) == ( 1'd1 )  ;
assign n2 =  ( n0 ) & ( n1 )  ;
assign n3 =  ( arg_0_TREADY ) == ( 1'd1 )  ;
assign n4 =  ( n2 ) & ( n3 )  ;
assign n5 =  ( arg_1_TREADY ) == ( 1'd0 )  ;
assign n6 =  ( arg_0_TREADY ) == ( 1'd0 )  ;
assign n7 =  ( n5 ) & ( n6 )  ;
assign n8 =  ( st_ready ) == ( 1'd0 )  ;
assign n9 =  ( n7 ) & ( n8 )  ;
assign n10 =  ( st_ready ) == ( 1'd1 )  ;
assign n11 =  ( n7 ) & ( n10 )  ;
assign n12 =  ( RAM_x ) == ( 9'd488 )  ;
assign n13 =  ( RAM_w ) == ( 3'd7 )  ;
assign n14 =  ( RAM_w ) + ( 3'd1 )  ;
assign n15 =  ( n13 ) ? ( 3'd0 ) : ( n14 ) ;
assign n16 =  ( n12 ) ? ( n15 ) : ( RAM_w ) ;
assign n17 =  ( arg_1_TVALID ) == ( 1'd1 )  ;
assign n18 =  ( arg_1_TREADY ) == ( 1'd1 )  ;
assign n19 =  ( n17 ) & ( n18 )  ;
assign n20 =  ( arg_0_TVALID ) == ( 1'd0 )  ;
assign n21 =  ( n19 ) & ( n20 )  ;
assign n22 =  ( n21 ) & ( n6 )  ;
assign n23 =  ( n22 ) ? ( RAM_w ) : ( RAM_w ) ;
assign n24 =  ( n11 ) ? ( n16 ) : ( n23 ) ;
assign n25 =  ( n9 ) ? ( RAM_w ) : ( n24 ) ;
assign n26 =  ( n4 ) ? ( RAM_w ) : ( n25 ) ;
assign n27 =  ( RAM_x ) == ( 9'd0 )  ;
assign n28 =  ( RAM_y ) == ( 10'd0 )  ;
assign n29 =  ( n27 ) & ( n28 )  ;
assign n30 =  ( RAM_x ) + ( 9'd1 )  ;
assign n31 =  ( n12 ) ? ( 9'd1 ) : ( n30 ) ;
assign n32 =  ( n29 ) ? ( 9'd1 ) : ( n31 ) ;
assign n33 =  ( n22 ) ? ( RAM_x ) : ( RAM_x ) ;
assign n34 =  ( n11 ) ? ( n32 ) : ( n33 ) ;
assign n35 =  ( n9 ) ? ( RAM_x ) : ( n34 ) ;
assign n36 =  ( n4 ) ? ( RAM_x ) : ( n35 ) ;
assign n37 =  ( RAM_y ) == ( 10'd648 )  ;
assign n38 =  ( RAM_y ) + ( 10'd1 )  ;
assign n39 =  ( n37 ) ? ( 10'd0 ) : ( n38 ) ;
assign n40 =  ( n12 ) ? ( n39 ) : ( RAM_y ) ;
assign n41 =  ( n22 ) ? ( RAM_y ) : ( RAM_y ) ;
assign n42 =  ( n11 ) ? ( n40 ) : ( n41 ) ;
assign n43 =  ( n9 ) ? ( RAM_y ) : ( n42 ) ;
assign n44 =  ( n4 ) ? ( RAM_y ) : ( n43 ) ;
assign n45 =  ( RAM_x ) == ( 9'd1 )  ;
assign n46 =  ( n45 ) & ( n37 )  ;
assign n47 =  ( RAM_x ) > ( 9'd8 )  ;
assign n48 =  ( RAM_y ) >= ( 10'd8 )  ;
assign n49 =  ( n47 ) & ( n48 )  ;
assign n50 =  ( RAM_y ) > ( 10'd8 )  ;
assign n51 =  ( n45 ) & ( n50 )  ;
assign n52 =  ( n49 ) | ( n51 )  ;
assign n53 = stencil_8[71:64] ;
assign n54 = stencil_7[71:64] ;
assign n55 = stencil_6[71:64] ;
assign n56 = stencil_5[71:64] ;
assign n57 = stencil_4[71:64] ;
assign n58 = stencil_3[71:64] ;
assign n59 = stencil_2[71:64] ;
assign n60 = stencil_1[71:64] ;
assign n61 = stencil_0[71:64] ;
assign n62 =  { ( n60 ) , ( n61 ) }  ;
assign n63 =  { ( n59 ) , ( n62 ) }  ;
assign n64 =  { ( n58 ) , ( n63 ) }  ;
assign n65 =  { ( n57 ) , ( n64 ) }  ;
assign n66 =  { ( n56 ) , ( n65 ) }  ;
assign n67 =  { ( n55 ) , ( n66 ) }  ;
assign n68 =  { ( n54 ) , ( n67 ) }  ;
assign n69 =  { ( n53 ) , ( n68 ) }  ;
assign n70 = stencil_8[63:56] ;
assign n71 = stencil_7[63:56] ;
assign n72 = stencil_6[63:56] ;
assign n73 = stencil_5[63:56] ;
assign n74 = stencil_4[63:56] ;
assign n75 = stencil_3[63:56] ;
assign n76 = stencil_2[63:56] ;
assign n77 = stencil_1[63:56] ;
assign n78 = stencil_0[63:56] ;
assign n79 =  { ( n77 ) , ( n78 ) }  ;
assign n80 =  { ( n76 ) , ( n79 ) }  ;
assign n81 =  { ( n75 ) , ( n80 ) }  ;
assign n82 =  { ( n74 ) , ( n81 ) }  ;
assign n83 =  { ( n73 ) , ( n82 ) }  ;
assign n84 =  { ( n72 ) , ( n83 ) }  ;
assign n85 =  { ( n71 ) , ( n84 ) }  ;
assign n86 =  { ( n70 ) , ( n85 ) }  ;
assign n87 = stencil_8[55:48] ;
assign n88 = stencil_7[55:48] ;
assign n89 = stencil_6[55:48] ;
assign n90 = stencil_5[55:48] ;
assign n91 = stencil_4[55:48] ;
assign n92 = stencil_3[55:48] ;
assign n93 = stencil_2[55:48] ;
assign n94 = stencil_1[55:48] ;
assign n95 = stencil_0[55:48] ;
assign n96 =  { ( n94 ) , ( n95 ) }  ;
assign n97 =  { ( n93 ) , ( n96 ) }  ;
assign n98 =  { ( n92 ) , ( n97 ) }  ;
assign n99 =  { ( n91 ) , ( n98 ) }  ;
assign n100 =  { ( n90 ) , ( n99 ) }  ;
assign n101 =  { ( n89 ) , ( n100 ) }  ;
assign n102 =  { ( n88 ) , ( n101 ) }  ;
assign n103 =  { ( n87 ) , ( n102 ) }  ;
assign n104 = stencil_8[47:40] ;
assign n105 = stencil_7[47:40] ;
assign n106 = stencil_6[47:40] ;
assign n107 = stencil_5[47:40] ;
assign n108 = stencil_4[47:40] ;
assign n109 = stencil_3[47:40] ;
assign n110 = stencil_2[47:40] ;
assign n111 = stencil_1[47:40] ;
assign n112 = stencil_0[47:40] ;
assign n113 =  { ( n111 ) , ( n112 ) }  ;
assign n114 =  { ( n110 ) , ( n113 ) }  ;
assign n115 =  { ( n109 ) , ( n114 ) }  ;
assign n116 =  { ( n108 ) , ( n115 ) }  ;
assign n117 =  { ( n107 ) , ( n116 ) }  ;
assign n118 =  { ( n106 ) , ( n117 ) }  ;
assign n119 =  { ( n105 ) , ( n118 ) }  ;
assign n120 =  { ( n104 ) , ( n119 ) }  ;
assign n121 = stencil_8[39:32] ;
assign n122 = stencil_7[39:32] ;
assign n123 = stencil_6[39:32] ;
assign n124 = stencil_5[39:32] ;
assign n125 = stencil_4[39:32] ;
assign n126 = stencil_3[39:32] ;
assign n127 = stencil_2[39:32] ;
assign n128 = stencil_1[39:32] ;
assign n129 = stencil_0[39:32] ;
assign n130 =  { ( n128 ) , ( n129 ) }  ;
assign n131 =  { ( n127 ) , ( n130 ) }  ;
assign n132 =  { ( n126 ) , ( n131 ) }  ;
assign n133 =  { ( n125 ) , ( n132 ) }  ;
assign n134 =  { ( n124 ) , ( n133 ) }  ;
assign n135 =  { ( n123 ) , ( n134 ) }  ;
assign n136 =  { ( n122 ) , ( n135 ) }  ;
assign n137 =  { ( n121 ) , ( n136 ) }  ;
assign n138 = stencil_8[31:24] ;
assign n139 = stencil_7[31:24] ;
assign n140 = stencil_6[31:24] ;
assign n141 = stencil_5[31:24] ;
assign n142 = stencil_4[31:24] ;
assign n143 = stencil_3[31:24] ;
assign n144 = stencil_2[31:24] ;
assign n145 = stencil_1[31:24] ;
assign n146 = stencil_0[31:24] ;
assign n147 =  { ( n145 ) , ( n146 ) }  ;
assign n148 =  { ( n144 ) , ( n147 ) }  ;
assign n149 =  { ( n143 ) , ( n148 ) }  ;
assign n150 =  { ( n142 ) , ( n149 ) }  ;
assign n151 =  { ( n141 ) , ( n150 ) }  ;
assign n152 =  { ( n140 ) , ( n151 ) }  ;
assign n153 =  { ( n139 ) , ( n152 ) }  ;
assign n154 =  { ( n138 ) , ( n153 ) }  ;
assign n155 = stencil_8[23:16] ;
assign n156 = stencil_7[23:16] ;
assign n157 = stencil_6[23:16] ;
assign n158 = stencil_5[23:16] ;
assign n159 = stencil_4[23:16] ;
assign n160 = stencil_3[23:16] ;
assign n161 = stencil_2[23:16] ;
assign n162 = stencil_1[23:16] ;
assign n163 = stencil_0[23:16] ;
assign n164 =  { ( n162 ) , ( n163 ) }  ;
assign n165 =  { ( n161 ) , ( n164 ) }  ;
assign n166 =  { ( n160 ) , ( n165 ) }  ;
assign n167 =  { ( n159 ) , ( n166 ) }  ;
assign n168 =  { ( n158 ) , ( n167 ) }  ;
assign n169 =  { ( n157 ) , ( n168 ) }  ;
assign n170 =  { ( n156 ) , ( n169 ) }  ;
assign n171 =  { ( n155 ) , ( n170 ) }  ;
assign n172 = stencil_8[15:8] ;
assign n173 = stencil_7[15:8] ;
assign n174 = stencil_6[15:8] ;
assign n175 = stencil_5[15:8] ;
assign n176 = stencil_4[15:8] ;
assign n177 = stencil_3[15:8] ;
assign n178 = stencil_2[15:8] ;
assign n179 = stencil_1[15:8] ;
assign n180 = stencil_0[15:8] ;
assign n181 =  { ( n179 ) , ( n180 ) }  ;
assign n182 =  { ( n178 ) , ( n181 ) }  ;
assign n183 =  { ( n177 ) , ( n182 ) }  ;
assign n184 =  { ( n176 ) , ( n183 ) }  ;
assign n185 =  { ( n175 ) , ( n184 ) }  ;
assign n186 =  { ( n174 ) , ( n185 ) }  ;
assign n187 =  { ( n173 ) , ( n186 ) }  ;
assign n188 =  { ( n172 ) , ( n187 ) }  ;
assign n189 = stencil_8[7:0] ;
assign n190 = stencil_7[7:0] ;
assign n191 = stencil_6[7:0] ;
assign n192 = stencil_5[7:0] ;
assign n193 = stencil_4[7:0] ;
assign n194 = stencil_3[7:0] ;
assign n195 = stencil_2[7:0] ;
assign n196 = stencil_1[7:0] ;
assign n197 = stencil_0[7:0] ;
assign n198 =  { ( n196 ) , ( n197 ) }  ;
assign n199 =  { ( n195 ) , ( n198 ) }  ;
assign n200 =  { ( n194 ) , ( n199 ) }  ;
assign n201 =  { ( n193 ) , ( n200 ) }  ;
assign n202 =  { ( n192 ) , ( n201 ) }  ;
assign n203 =  { ( n191 ) , ( n202 ) }  ;
assign n204 =  { ( n190 ) , ( n203 ) }  ;
assign n205 =  { ( n189 ) , ( n204 ) }  ;
assign n206 =  { ( n188 ) , ( n205 ) }  ;
assign n207 =  { ( n171 ) , ( n206 ) }  ;
assign n208 =  { ( n154 ) , ( n207 ) }  ;
assign n209 =  { ( n137 ) , ( n208 ) }  ;
assign n210 =  { ( n120 ) , ( n209 ) }  ;
assign n211 =  { ( n103 ) , ( n210 ) }  ;
assign n212 =  { ( n86 ) , ( n211 ) }  ;
assign n213 =  { ( n69 ) , ( n212 ) }  ;
assign n214 =  ( n52 ) ? ( n213 ) : ( proc_in ) ;
assign n215 =  ( n46 ) ? ( proc_in ) : ( n214 ) ;
fun_gb_fun  applyFunc_n217(
    .arg1( n215 ),
    .result( n216 )
);
assign n218 = n216 ;
assign n219 =  ( n46 ) ? ( arg_0_TDATA ) : ( n218 ) ;
assign n220 =  ( n22 ) ? ( arg_0_TDATA ) : ( arg_0_TDATA ) ;
assign n221 =  ( n11 ) ? ( arg_0_TDATA ) : ( n220 ) ;
assign n222 =  ( n9 ) ? ( n219 ) : ( n221 ) ;
assign n223 =  ( n4 ) ? ( arg_0_TDATA ) : ( n222 ) ;
assign n224 =  ( gbit ) == ( 4'd0 )  ;
assign n225 =  ( gbit ) == ( 4'd7 )  ;
assign n226 =  ( n224 ) | ( n225 )  ;
assign n227 =  ( n226 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n228 =  ( n52 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n229 =  ( n46 ) ? ( arg_0_TVALID ) : ( n228 ) ;
assign n230 =  ( n29 ) ? ( 1'd0 ) : ( arg_0_TVALID ) ;
assign n231 =  ( n22 ) ? ( 1'd0 ) : ( arg_0_TVALID ) ;
assign n232 =  ( n11 ) ? ( n230 ) : ( n231 ) ;
assign n233 =  ( n9 ) ? ( n229 ) : ( n232 ) ;
assign n234 =  ( n4 ) ? ( n227 ) : ( n233 ) ;
assign n235 =  ( 9'd488 ) - ( 9'd1 )  ;
assign n236 =  ( RAM_x ) == ( n235 )  ;
assign n237 =  ( 10'd648 ) - ( 10'd1 )  ;
assign n238 =  ( RAM_y ) == ( n237 )  ;
assign n239 =  ( n236 ) & ( n238 )  ;
assign n240 =  ( n239 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n241 =  ( RAM_y ) < ( 10'd8 )  ;
assign n242 =  ( n241 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n243 =  ( n29 ) ? ( 1'd1 ) : ( n242 ) ;
assign n244 =  ( n22 ) ? ( 1'd0 ) : ( arg_1_TREADY ) ;
assign n245 =  ( n11 ) ? ( n243 ) : ( n244 ) ;
assign n246 =  ( n9 ) ? ( n240 ) : ( n245 ) ;
assign n247 =  ( n4 ) ? ( arg_1_TREADY ) : ( n246 ) ;
assign n248 =  ( n22 ) ? ( arg_1_TDATA ) : ( cur_pix ) ;
assign n249 =  ( n11 ) ? ( cur_pix ) : ( n248 ) ;
assign n250 =  ( n9 ) ? ( cur_pix ) : ( n249 ) ;
assign n251 =  ( n4 ) ? ( cur_pix ) : ( n250 ) ;
assign n252 =  ( n12 ) & ( n37 )  ;
assign n253 =  ( gbit ) + ( 4'd1 )  ;
assign n254 =  ( n252 ) ? ( n253 ) : ( gbit ) ;
assign n255 =  ( n4 ) ? ( n254 ) : ( gbit ) ;
assign n256 =  ( n11 ) ? ( cur_pix ) : ( pre_pix ) ;
assign n257 =  ( n9 ) ? ( pre_pix ) : ( n256 ) ;
assign n258 =  ( n11 ) ? ( proc_in ) : ( proc_in ) ;
assign n259 =  ( n9 ) ? ( n215 ) : ( n258 ) ;
assign n260 =  ( n11 ) ? ( n243 ) : ( st_ready ) ;
assign n261 =  ( n9 ) ? ( 1'd1 ) : ( n260 ) ;
assign n262 =  ( n241 ) ? ( stencil_0 ) : ( stencil_1 ) ;
assign n263 =  ( n22 ) ? ( stencil_0 ) : ( stencil_0 ) ;
assign n264 =  ( n11 ) ? ( stencil_0 ) : ( n263 ) ;
assign n265 =  ( n9 ) ? ( n262 ) : ( n264 ) ;
assign n266 =  ( n4 ) ? ( stencil_0 ) : ( n265 ) ;
assign n267 =  ( n241 ) ? ( stencil_1 ) : ( stencil_2 ) ;
assign n268 =  ( n22 ) ? ( stencil_1 ) : ( stencil_1 ) ;
assign n269 =  ( n11 ) ? ( stencil_1 ) : ( n268 ) ;
assign n270 =  ( n9 ) ? ( n267 ) : ( n269 ) ;
assign n271 =  ( n4 ) ? ( stencil_1 ) : ( n270 ) ;
assign n272 =  ( n241 ) ? ( stencil_2 ) : ( stencil_3 ) ;
assign n273 =  ( n22 ) ? ( stencil_2 ) : ( stencil_2 ) ;
assign n274 =  ( n11 ) ? ( stencil_2 ) : ( n273 ) ;
assign n275 =  ( n9 ) ? ( n272 ) : ( n274 ) ;
assign n276 =  ( n4 ) ? ( stencil_2 ) : ( n275 ) ;
assign n277 =  ( n241 ) ? ( stencil_3 ) : ( stencil_4 ) ;
assign n278 =  ( n22 ) ? ( stencil_3 ) : ( stencil_3 ) ;
assign n279 =  ( n11 ) ? ( stencil_3 ) : ( n278 ) ;
assign n280 =  ( n9 ) ? ( n277 ) : ( n279 ) ;
assign n281 =  ( n4 ) ? ( stencil_3 ) : ( n280 ) ;
assign n282 =  ( n241 ) ? ( stencil_4 ) : ( stencil_5 ) ;
assign n283 =  ( n22 ) ? ( stencil_4 ) : ( stencil_4 ) ;
assign n284 =  ( n11 ) ? ( stencil_4 ) : ( n283 ) ;
assign n285 =  ( n9 ) ? ( n282 ) : ( n284 ) ;
assign n286 =  ( n4 ) ? ( stencil_4 ) : ( n285 ) ;
assign n287 =  ( n241 ) ? ( stencil_5 ) : ( stencil_6 ) ;
assign n288 =  ( n22 ) ? ( stencil_5 ) : ( stencil_5 ) ;
assign n289 =  ( n11 ) ? ( stencil_5 ) : ( n288 ) ;
assign n290 =  ( n9 ) ? ( n287 ) : ( n289 ) ;
assign n291 =  ( n4 ) ? ( stencil_5 ) : ( n290 ) ;
assign n292 =  ( n241 ) ? ( stencil_6 ) : ( stencil_7 ) ;
assign n293 =  ( n22 ) ? ( stencil_6 ) : ( stencil_6 ) ;
assign n294 =  ( n11 ) ? ( stencil_6 ) : ( n293 ) ;
assign n295 =  ( n9 ) ? ( n292 ) : ( n294 ) ;
assign n296 =  ( n4 ) ? ( stencil_6 ) : ( n295 ) ;
assign n297 =  ( n241 ) ? ( stencil_7 ) : ( stencil_8 ) ;
assign n298 =  ( n22 ) ? ( stencil_7 ) : ( stencil_7 ) ;
assign n299 =  ( n11 ) ? ( stencil_7 ) : ( n298 ) ;
assign n300 =  ( n9 ) ? ( n297 ) : ( n299 ) ;
assign n301 =  ( n4 ) ? ( stencil_7 ) : ( n300 ) ;
assign n302 =  ( RAM_w ) == ( 3'd0 )  ;
assign n303 =  ( RAM_x ) - ( 9'd1 )  ;
assign n304 =  (  RAM_7 [ n303 ] )  ;
assign n305 =  ( RAM_w ) == ( 3'd1 )  ;
assign n306 =  (  RAM_0 [ n303 ] )  ;
assign n307 =  ( RAM_w ) == ( 3'd2 )  ;
assign n308 =  (  RAM_1 [ n303 ] )  ;
assign n309 =  ( RAM_w ) == ( 3'd3 )  ;
assign n310 =  (  RAM_2 [ n303 ] )  ;
assign n311 =  ( RAM_w ) == ( 3'd4 )  ;
assign n312 =  (  RAM_3 [ n303 ] )  ;
assign n313 =  ( RAM_w ) == ( 3'd5 )  ;
assign n314 =  (  RAM_4 [ n303 ] )  ;
assign n315 =  ( RAM_w ) == ( 3'd6 )  ;
assign n316 =  (  RAM_5 [ n303 ] )  ;
assign n317 =  (  RAM_6 [ n303 ] )  ;
assign n318 =  ( n315 ) ? ( n316 ) : ( n317 ) ;
assign n319 =  ( n313 ) ? ( n314 ) : ( n318 ) ;
assign n320 =  ( n311 ) ? ( n312 ) : ( n319 ) ;
assign n321 =  ( n309 ) ? ( n310 ) : ( n320 ) ;
assign n322 =  ( n307 ) ? ( n308 ) : ( n321 ) ;
assign n323 =  ( n305 ) ? ( n306 ) : ( n322 ) ;
assign n324 =  ( n302 ) ? ( n304 ) : ( n323 ) ;
assign n325 =  ( n315 ) ? ( n314 ) : ( n316 ) ;
assign n326 =  ( n313 ) ? ( n312 ) : ( n325 ) ;
assign n327 =  ( n311 ) ? ( n310 ) : ( n326 ) ;
assign n328 =  ( n309 ) ? ( n308 ) : ( n327 ) ;
assign n329 =  ( n307 ) ? ( n306 ) : ( n328 ) ;
assign n330 =  ( n305 ) ? ( n304 ) : ( n329 ) ;
assign n331 =  ( n302 ) ? ( n317 ) : ( n330 ) ;
assign n332 =  ( n315 ) ? ( n312 ) : ( n314 ) ;
assign n333 =  ( n313 ) ? ( n310 ) : ( n332 ) ;
assign n334 =  ( n311 ) ? ( n308 ) : ( n333 ) ;
assign n335 =  ( n309 ) ? ( n306 ) : ( n334 ) ;
assign n336 =  ( n307 ) ? ( n304 ) : ( n335 ) ;
assign n337 =  ( n305 ) ? ( n317 ) : ( n336 ) ;
assign n338 =  ( n302 ) ? ( n316 ) : ( n337 ) ;
assign n339 =  ( n315 ) ? ( n310 ) : ( n312 ) ;
assign n340 =  ( n313 ) ? ( n308 ) : ( n339 ) ;
assign n341 =  ( n311 ) ? ( n306 ) : ( n340 ) ;
assign n342 =  ( n309 ) ? ( n304 ) : ( n341 ) ;
assign n343 =  ( n307 ) ? ( n317 ) : ( n342 ) ;
assign n344 =  ( n305 ) ? ( n316 ) : ( n343 ) ;
assign n345 =  ( n302 ) ? ( n314 ) : ( n344 ) ;
assign n346 =  ( n315 ) ? ( n308 ) : ( n310 ) ;
assign n347 =  ( n313 ) ? ( n306 ) : ( n346 ) ;
assign n348 =  ( n311 ) ? ( n304 ) : ( n347 ) ;
assign n349 =  ( n309 ) ? ( n317 ) : ( n348 ) ;
assign n350 =  ( n307 ) ? ( n316 ) : ( n349 ) ;
assign n351 =  ( n305 ) ? ( n314 ) : ( n350 ) ;
assign n352 =  ( n302 ) ? ( n312 ) : ( n351 ) ;
assign n353 =  ( n315 ) ? ( n306 ) : ( n308 ) ;
assign n354 =  ( n313 ) ? ( n304 ) : ( n353 ) ;
assign n355 =  ( n311 ) ? ( n317 ) : ( n354 ) ;
assign n356 =  ( n309 ) ? ( n316 ) : ( n355 ) ;
assign n357 =  ( n307 ) ? ( n314 ) : ( n356 ) ;
assign n358 =  ( n305 ) ? ( n312 ) : ( n357 ) ;
assign n359 =  ( n302 ) ? ( n310 ) : ( n358 ) ;
assign n360 =  ( n315 ) ? ( n304 ) : ( n306 ) ;
assign n361 =  ( n313 ) ? ( n317 ) : ( n360 ) ;
assign n362 =  ( n311 ) ? ( n316 ) : ( n361 ) ;
assign n363 =  ( n309 ) ? ( n314 ) : ( n362 ) ;
assign n364 =  ( n307 ) ? ( n312 ) : ( n363 ) ;
assign n365 =  ( n305 ) ? ( n310 ) : ( n364 ) ;
assign n366 =  ( n302 ) ? ( n308 ) : ( n365 ) ;
assign n367 =  ( n315 ) ? ( n317 ) : ( n304 ) ;
assign n368 =  ( n313 ) ? ( n316 ) : ( n367 ) ;
assign n369 =  ( n311 ) ? ( n314 ) : ( n368 ) ;
assign n370 =  ( n309 ) ? ( n312 ) : ( n369 ) ;
assign n371 =  ( n307 ) ? ( n310 ) : ( n370 ) ;
assign n372 =  ( n305 ) ? ( n308 ) : ( n371 ) ;
assign n373 =  ( n302 ) ? ( n306 ) : ( n372 ) ;
assign n374 =  { ( n366 ) , ( n373 ) }  ;
assign n375 =  { ( n359 ) , ( n374 ) }  ;
assign n376 =  { ( n352 ) , ( n375 ) }  ;
assign n377 =  { ( n345 ) , ( n376 ) }  ;
assign n378 =  { ( n338 ) , ( n377 ) }  ;
assign n379 =  { ( n331 ) , ( n378 ) }  ;
assign n380 =  { ( n324 ) , ( n379 ) }  ;
assign n381 =  { ( pre_pix ) , ( n380 ) }  ;
assign n382 =  ( n241 ) ? ( stencil_8 ) : ( n381 ) ;
assign n383 =  ( n22 ) ? ( stencil_8 ) : ( stencil_8 ) ;
assign n384 =  ( n11 ) ? ( n382 ) : ( n383 ) ;
assign n385 =  ( n9 ) ? ( stencil_8 ) : ( n384 ) ;
assign n386 =  ( n4 ) ? ( stencil_8 ) : ( n385 ) ;
assign n387 = ~ ( n4 ) ;
assign n388 =  ( 1'b1 ) & ( n387 )  ;
assign n389 = ~ ( n9 ) ;
assign n390 =  ( n388 ) & ( n389 )  ;
assign n391 = ~ ( n11 ) ;
assign n392 =  ( n390 ) & ( n391 )  ;
assign n393 = ~ ( n22 ) ;
assign n394 =  ( n392 ) & ( n393 )  ;
assign n395 =  ( n392 ) & ( n22 )  ;
assign n396 =  ( n390 ) & ( n11 )  ;
assign n397 = ~ ( n29 ) ;
assign n398 =  ( n396 ) & ( n397 )  ;
assign n399 = ~ ( n302 ) ;
assign n400 =  ( n398 ) & ( n399 )  ;
assign n401 =  ( n398 ) & ( n302 )  ;
assign n402 =  ( n396 ) & ( n29 )  ;
assign n403 =  ( n388 ) & ( n9 )  ;
assign n404 =  ( 1'b1 ) & ( n4 )  ;
assign RAM_0_addr0 = n401 ? (n303) : (0);
assign RAM_0_data0 = n401 ? (pre_pix) : ('dx);
assign RAM_0_wen0 = n401 ? ( 1'b1 ) : (1'b0);
assign n405 = ~ ( n305 ) ;
assign n406 =  ( n398 ) & ( n405 )  ;
assign n407 =  ( n398 ) & ( n305 )  ;
assign RAM_1_addr0 = n407 ? (n303) : (0);
assign RAM_1_data0 = n407 ? (pre_pix) : ('dx);
assign RAM_1_wen0 = n407 ? ( 1'b1 ) : (1'b0);
assign n408 = ~ ( n307 ) ;
assign n409 =  ( n398 ) & ( n408 )  ;
assign n410 =  ( n398 ) & ( n307 )  ;
assign RAM_2_addr0 = n410 ? (n303) : (0);
assign RAM_2_data0 = n410 ? (pre_pix) : ('dx);
assign RAM_2_wen0 = n410 ? ( 1'b1 ) : (1'b0);
assign n411 = ~ ( n309 ) ;
assign n412 =  ( n398 ) & ( n411 )  ;
assign n413 =  ( n398 ) & ( n309 )  ;
assign RAM_3_addr0 = n413 ? (n303) : (0);
assign RAM_3_data0 = n413 ? (pre_pix) : ('dx);
assign RAM_3_wen0 = n413 ? ( 1'b1 ) : (1'b0);
assign n414 = ~ ( n311 ) ;
assign n415 =  ( n398 ) & ( n414 )  ;
assign n416 =  ( n398 ) & ( n311 )  ;
assign RAM_4_addr0 = n416 ? (n303) : (0);
assign RAM_4_data0 = n416 ? (pre_pix) : ('dx);
assign RAM_4_wen0 = n416 ? ( 1'b1 ) : (1'b0);
assign n417 = ~ ( n313 ) ;
assign n418 =  ( n398 ) & ( n417 )  ;
assign n419 =  ( n398 ) & ( n313 )  ;
assign RAM_5_addr0 = n419 ? (n303) : (0);
assign RAM_5_data0 = n419 ? (pre_pix) : ('dx);
assign RAM_5_wen0 = n419 ? ( 1'b1 ) : (1'b0);
assign n420 = ~ ( n315 ) ;
assign n421 =  ( n398 ) & ( n420 )  ;
assign n422 =  ( n398 ) & ( n315 )  ;
assign RAM_6_addr0 = n422 ? (n303) : (0);
assign RAM_6_data0 = n422 ? (pre_pix) : ('dx);
assign RAM_6_wen0 = n422 ? ( 1'b1 ) : (1'b0);
assign n423 = ~ ( n13 ) ;
assign n424 =  ( n398 ) & ( n423 )  ;
assign n425 =  ( n398 ) & ( n13 )  ;
assign RAM_7_addr0 = n425 ? (n303) : (0);
assign RAM_7_data0 = n425 ? (pre_pix) : ('dx);
assign RAM_7_wen0 = n425 ? ( 1'b1 ) : (1'b0);
always @(posedge clk) begin
   if(rst) begin
       RAM_w <= RAM_w;
       RAM_x <= RAM_x;
       RAM_y <= RAM_y;
       arg_0_TDATA <= arg_0_TDATA;
       arg_0_TVALID <= arg_0_TVALID;
       arg_1_TREADY <= arg_1_TREADY;
       cur_pix <= cur_pix;
       gbit <= gbit;
       pre_pix <= pre_pix;
       proc_in <= proc_in;
       st_ready <= st_ready;
       stencil_0 <= stencil_0;
       stencil_1 <= stencil_1;
       stencil_2 <= stencil_2;
       stencil_3 <= stencil_3;
       stencil_4 <= stencil_4;
       stencil_5 <= stencil_5;
       stencil_6 <= stencil_6;
       stencil_7 <= stencil_7;
       stencil_8 <= stencil_8;
   end
   else if(step) begin
       RAM_w <= n26;
       RAM_x <= n36;
       RAM_y <= n44;
       arg_0_TDATA <= n223;
       arg_0_TVALID <= n234;
       arg_1_TREADY <= n247;
       cur_pix <= n251;
       gbit <= n255;
       pre_pix <= n257;
       proc_in <= n259;
       st_ready <= n261;
       stencil_0 <= n266;
       stencil_1 <= n271;
       stencil_2 <= n276;
       stencil_3 <= n281;
       stencil_4 <= n286;
       stencil_5 <= n291;
       stencil_6 <= n296;
       stencil_7 <= n301;
       stencil_8 <= n386;
       if (RAM_0_wen0) begin
           RAM_0 [ RAM_0_addr0 ] <= RAM_0_data0 ;
       end
       if (RAM_1_wen0) begin
           RAM_1 [ RAM_1_addr0 ] <= RAM_1_data0 ;
       end
       if (RAM_2_wen0) begin
           RAM_2 [ RAM_2_addr0 ] <= RAM_2_data0 ;
       end
       if (RAM_3_wen0) begin
           RAM_3 [ RAM_3_addr0 ] <= RAM_3_data0 ;
       end
       if (RAM_4_wen0) begin
           RAM_4 [ RAM_4_addr0 ] <= RAM_4_data0 ;
       end
       if (RAM_5_wen0) begin
           RAM_5 [ RAM_5_addr0 ] <= RAM_5_data0 ;
       end
       if (RAM_6_wen0) begin
           RAM_6 [ RAM_6_addr0 ] <= RAM_6_data0 ;
       end
       if (RAM_7_wen0) begin
           RAM_7 [ RAM_7_addr0 ] <= RAM_7_data0 ;
       end
   end
end
endmodule
