module SPEC_B(
arg_0_TREADY,
arg_1_TDATA,
arg_1_TVALID,
LB1D_buff,
LB1D_in,
LB1D_it_1,
LB1D_p_cnt,
LB1D_uIn,
LB2D_proc_w,
LB2D_proc_x,
LB2D_proc_y,
LB2D_shift_0,
LB2D_shift_1,
LB2D_shift_2,
LB2D_shift_3,
LB2D_shift_4,
LB2D_shift_5,
LB2D_shift_6,
LB2D_shift_7,
LB2D_shift_x,
LB2D_shift_y,
arg_0_TDATA,
arg_0_TVALID,
arg_1_TREADY,
gb_exit_it_1,
gb_exit_it_2,
gb_exit_it_3,
gb_exit_it_4,
gb_exit_it_5,
gb_exit_it_6,
gb_exit_it_7,
gb_exit_it_8,
gb_p_cnt,
gb_pp_it_1,
gb_pp_it_2,
gb_pp_it_3,
gb_pp_it_4,
gb_pp_it_5,
gb_pp_it_6,
gb_pp_it_7,
gb_pp_it_8,
gb_pp_it_9,
in_stream_buff_0,
in_stream_buff_1,
in_stream_empty,
in_stream_full,
slice_stream_buff_0,
slice_stream_buff_1,
slice_stream_empty,
slice_stream_full,
stencil_stream_buff_0,
stencil_stream_buff_1,
stencil_stream_empty,
stencil_stream_full,
clk,rst,
step
);
input            arg_0_TREADY;
input      [7:0] arg_1_TDATA;
input            arg_1_TVALID;
input clk;
input rst;
input step;
output      [7:0] LB1D_buff;
output      [7:0] LB1D_in;
output            LB1D_it_1;
output     [18:0] LB1D_p_cnt;
output      [7:0] LB1D_uIn;
output     [63:0] LB2D_proc_w;
output      [8:0] LB2D_proc_x;
output      [9:0] LB2D_proc_y;
output     [71:0] LB2D_shift_0;
output     [71:0] LB2D_shift_1;
output     [71:0] LB2D_shift_2;
output     [71:0] LB2D_shift_3;
output     [71:0] LB2D_shift_4;
output     [71:0] LB2D_shift_5;
output     [71:0] LB2D_shift_6;
output     [71:0] LB2D_shift_7;
output      [8:0] LB2D_shift_x;
output      [9:0] LB2D_shift_y;
output      [7:0] arg_0_TDATA;
output            arg_0_TVALID;
output            arg_1_TREADY;
output            gb_exit_it_1;
output            gb_exit_it_2;
output            gb_exit_it_3;
output            gb_exit_it_4;
output            gb_exit_it_5;
output            gb_exit_it_6;
output            gb_exit_it_7;
output            gb_exit_it_8;
output     [18:0] gb_p_cnt;
output            gb_pp_it_1;
output            gb_pp_it_2;
output            gb_pp_it_3;
output            gb_pp_it_4;
output            gb_pp_it_5;
output            gb_pp_it_6;
output            gb_pp_it_7;
output            gb_pp_it_8;
output            gb_pp_it_9;
output      [7:0] in_stream_buff_0;
output      [7:0] in_stream_buff_1;
output            in_stream_empty;
output            in_stream_full;
output     [71:0] slice_stream_buff_0;
output     [71:0] slice_stream_buff_1;
output            slice_stream_empty;
output            slice_stream_full;
output    [647:0] stencil_stream_buff_0;
output    [647:0] stencil_stream_buff_1;
output            stencil_stream_empty;
output            stencil_stream_full;
reg      [7:0] LB1D_buff;
reg      [7:0] LB1D_in;
reg            LB1D_it_1;
reg     [18:0] LB1D_p_cnt;
reg      [7:0] LB1D_uIn;
reg     [63:0] LB2D_proc_w;
reg      [8:0] LB2D_proc_x;
reg      [9:0] LB2D_proc_y;
reg     [71:0] LB2D_shift_0;
reg     [71:0] LB2D_shift_1;
reg     [71:0] LB2D_shift_2;
reg     [71:0] LB2D_shift_3;
reg     [71:0] LB2D_shift_4;
reg     [71:0] LB2D_shift_5;
reg     [71:0] LB2D_shift_6;
reg     [71:0] LB2D_shift_7;
reg      [8:0] LB2D_shift_x;
reg      [9:0] LB2D_shift_y;
reg      [7:0] arg_0_TDATA;
reg            arg_0_TVALID;
reg            arg_1_TREADY;
reg            gb_exit_it_1;
reg            gb_exit_it_2;
reg            gb_exit_it_3;
reg            gb_exit_it_4;
reg            gb_exit_it_5;
reg            gb_exit_it_6;
reg            gb_exit_it_7;
reg            gb_exit_it_8;
reg     [18:0] gb_p_cnt;
reg            gb_pp_it_1;
reg            gb_pp_it_2;
reg            gb_pp_it_3;
reg            gb_pp_it_4;
reg            gb_pp_it_5;
reg            gb_pp_it_6;
reg            gb_pp_it_7;
reg            gb_pp_it_8;
reg            gb_pp_it_9;
reg      [7:0] in_stream_buff_0;
reg      [7:0] in_stream_buff_1;
reg            in_stream_empty;
reg            in_stream_full;
reg     [71:0] slice_stream_buff_0;
reg     [71:0] slice_stream_buff_1;
reg            slice_stream_empty;
reg            slice_stream_full;
reg    [647:0] stencil_stream_buff_0;
reg    [647:0] stencil_stream_buff_1;
reg            stencil_stream_empty;
reg            stencil_stream_full;
wire            arg_0_TREADY;
wire      [7:0] arg_1_TDATA;
wire            arg_1_TVALID;
wire            n0;
wire            n1;
wire            n2;
wire            n3;
wire            n4;
wire            n5;
wire            n6;
wire            n7;
wire            n8;
wire            n9;
wire            n10;
wire            n11;
wire            n12;
wire            n13;
wire            n14;
wire            n15;
wire            n16;
wire            n17;
wire            n18;
wire            n19;
wire            n20;
wire            n21;
wire            n22;
wire            n23;
wire            n24;
wire            n25;
wire            n26;
wire            n27;
wire            n28;
wire            n29;
wire            n30;
wire            n31;
wire            n32;
wire            n33;
wire            n34;
wire            n35;
wire            n36;
wire            n37;
wire            n38;
wire            n39;
wire            n40;
wire            n41;
wire            n42;
wire            n43;
wire      [7:0] n44;
wire      [7:0] n45;
wire      [7:0] n46;
wire      [7:0] n47;
wire      [7:0] n48;
wire      [7:0] n49;
wire      [7:0] n50;
wire      [7:0] n51;
wire      [7:0] n52;
wire      [7:0] n53;
wire      [7:0] n54;
wire      [7:0] n55;
wire      [7:0] n56;
wire      [7:0] n57;
wire      [7:0] n58;
wire      [7:0] n59;
wire            n60;
wire            n61;
wire            n62;
wire     [18:0] n63;
wire     [18:0] n64;
wire     [18:0] n65;
wire     [18:0] n66;
wire     [18:0] n67;
wire     [18:0] n68;
wire     [18:0] n69;
wire     [18:0] n70;
wire     [18:0] n71;
wire      [7:0] n72;
wire      [7:0] n73;
wire      [7:0] n74;
wire      [7:0] n75;
wire      [7:0] n76;
wire      [7:0] n77;
wire      [7:0] n78;
wire            n79;
wire            n80;
wire     [63:0] n81;
wire     [63:0] n82;
wire     [63:0] n83;
wire     [63:0] n84;
wire     [63:0] n85;
wire     [63:0] n86;
wire     [63:0] n87;
wire     [63:0] n88;
wire     [63:0] n89;
wire     [63:0] n90;
wire      [8:0] n91;
wire      [8:0] n92;
wire      [8:0] n93;
wire      [8:0] n94;
wire      [8:0] n95;
wire      [8:0] n96;
wire      [8:0] n97;
wire      [8:0] n98;
wire      [8:0] n99;
wire            n100;
wire      [9:0] n101;
wire      [9:0] n102;
wire      [9:0] n103;
wire      [9:0] n104;
wire      [9:0] n105;
wire      [9:0] n106;
wire      [9:0] n107;
wire      [9:0] n108;
wire      [9:0] n109;
wire      [9:0] n110;
wire     [71:0] n111;
wire     [71:0] n112;
wire     [71:0] n113;
wire     [71:0] n114;
wire     [71:0] n115;
wire     [71:0] n116;
wire     [71:0] n117;
wire     [71:0] n118;
wire     [71:0] n119;
wire     [71:0] n120;
wire     [71:0] n121;
wire     [71:0] n122;
wire     [71:0] n123;
wire     [71:0] n124;
wire     [71:0] n125;
wire     [71:0] n126;
wire     [71:0] n127;
wire     [71:0] n128;
wire     [71:0] n129;
wire     [71:0] n130;
wire     [71:0] n131;
wire     [71:0] n132;
wire     [71:0] n133;
wire     [71:0] n134;
wire     [71:0] n135;
wire     [71:0] n136;
wire     [71:0] n137;
wire     [71:0] n138;
wire     [71:0] n139;
wire     [71:0] n140;
wire     [71:0] n141;
wire     [71:0] n142;
wire     [71:0] n143;
wire     [71:0] n144;
wire     [71:0] n145;
wire     [71:0] n146;
wire     [71:0] n147;
wire     [71:0] n148;
wire     [71:0] n149;
wire     [71:0] n150;
wire     [71:0] n151;
wire     [71:0] n152;
wire     [71:0] n153;
wire     [71:0] n154;
wire     [71:0] n155;
wire     [71:0] n156;
wire     [71:0] n157;
wire     [71:0] n158;
wire     [71:0] n159;
wire            n160;
wire     [71:0] n161;
wire     [71:0] n162;
wire     [71:0] n163;
wire     [71:0] n164;
wire     [71:0] n165;
wire     [71:0] n166;
wire     [71:0] n167;
wire     [71:0] n168;
wire            n169;
wire            n170;
wire            n171;
wire            n172;
wire      [8:0] n173;
wire      [8:0] n174;
wire      [8:0] n175;
wire      [8:0] n176;
wire      [8:0] n177;
wire      [8:0] n178;
wire      [8:0] n179;
wire      [8:0] n180;
wire      [8:0] n181;
wire            n182;
wire            n183;
wire      [9:0] n184;
wire      [9:0] n185;
wire      [9:0] n186;
wire      [9:0] n187;
wire      [9:0] n188;
wire      [9:0] n189;
wire      [9:0] n190;
wire      [9:0] n191;
wire      [9:0] n192;
wire      [9:0] n193;
wire            n194;
wire    [647:0] n195;
wire      [7:0] n196;
wire      [7:0] n197;
wire      [7:0] n198;
wire      [7:0] n199;
wire      [7:0] n200;
wire      [7:0] n201;
wire      [7:0] n202;
wire      [7:0] n203;
wire            n204;
wire            n205;
wire            n206;
wire            n207;
wire            n208;
wire            n209;
wire            n210;
wire            n211;
wire            n212;
wire            n213;
wire            n214;
wire            n215;
wire            n216;
wire            n217;
wire            n218;
wire            n219;
wire            n220;
wire            n221;
wire            n222;
wire            n223;
wire            n224;
wire            n225;
wire            n226;
wire            n227;
wire            n228;
wire            n229;
wire            n230;
wire            n231;
wire            n232;
wire            n233;
wire            n234;
wire            n235;
wire            n236;
wire            n237;
wire            n238;
wire            n239;
wire            n240;
wire            n241;
wire            n242;
wire            n243;
wire            n244;
wire            n245;
wire            n246;
wire            n247;
wire            n248;
wire            n249;
wire            n250;
wire            n251;
wire            n252;
wire            n253;
wire            n254;
wire            n255;
wire            n256;
wire            n257;
wire            n258;
wire            n259;
wire            n260;
wire            n261;
wire            n262;
wire            n263;
wire            n264;
wire            n265;
wire            n266;
wire            n267;
wire            n268;
wire            n269;
wire            n270;
wire            n271;
wire            n272;
wire            n273;
wire            n274;
wire            n275;
wire            n276;
wire            n277;
wire            n278;
wire            n279;
wire            n280;
wire            n281;
wire     [18:0] n282;
wire     [18:0] n283;
wire     [18:0] n284;
wire     [18:0] n285;
wire     [18:0] n286;
wire     [18:0] n287;
wire     [18:0] n288;
wire     [18:0] n289;
wire     [18:0] n290;
wire            n291;
wire            n292;
wire            n293;
wire            n294;
wire            n295;
wire            n296;
wire            n297;
wire            n298;
wire            n299;
wire            n300;
wire            n301;
wire            n302;
wire            n303;
wire            n304;
wire            n305;
wire            n306;
wire            n307;
wire            n308;
wire            n309;
wire            n310;
wire            n311;
wire            n312;
wire            n313;
wire            n314;
wire            n315;
wire            n316;
wire            n317;
wire            n318;
wire            n319;
wire            n320;
wire            n321;
wire            n322;
wire            n323;
wire            n324;
wire            n325;
wire            n326;
wire            n327;
wire            n328;
wire            n329;
wire            n330;
wire            n331;
wire            n332;
wire            n333;
wire            n334;
wire            n335;
wire            n336;
wire            n337;
wire            n338;
wire            n339;
wire            n340;
wire            n341;
wire            n342;
wire            n343;
wire            n344;
wire            n345;
wire            n346;
wire            n347;
wire            n348;
wire            n349;
wire            n350;
wire            n351;
wire            n352;
wire            n353;
wire      [7:0] n354;
wire      [7:0] n355;
wire      [7:0] n356;
wire      [7:0] n357;
wire      [7:0] n358;
wire      [7:0] n359;
wire      [7:0] n360;
wire      [7:0] n361;
wire      [7:0] n362;
wire      [7:0] n363;
wire      [7:0] n364;
wire      [7:0] n365;
wire      [7:0] n366;
wire      [7:0] n367;
wire            n368;
wire            n369;
wire            n370;
wire            n371;
wire            n372;
wire            n373;
wire            n374;
wire            n375;
wire            n376;
wire            n377;
wire            n378;
wire            n379;
wire            n380;
wire            n381;
wire            n382;
wire            n383;
wire            n384;
wire            n385;
wire      [7:0] n386;
wire            n387;
wire      [8:0] n388;
wire      [7:0] n389;
wire            n390;
wire      [7:0] n391;
wire            n392;
wire      [7:0] n393;
wire            n394;
wire      [7:0] n395;
wire            n396;
wire      [7:0] n397;
wire            n398;
wire      [7:0] n399;
wire            n400;
wire      [7:0] n401;
wire      [7:0] n402;
wire      [7:0] n403;
wire      [7:0] n404;
wire      [7:0] n405;
wire      [7:0] n406;
wire      [7:0] n407;
wire      [7:0] n408;
wire      [7:0] n409;
wire      [7:0] n410;
wire      [7:0] n411;
wire      [7:0] n412;
wire      [7:0] n413;
wire      [7:0] n414;
wire      [7:0] n415;
wire      [7:0] n416;
wire      [7:0] n417;
wire      [7:0] n418;
wire      [7:0] n419;
wire      [7:0] n420;
wire      [7:0] n421;
wire      [7:0] n422;
wire      [7:0] n423;
wire      [7:0] n424;
wire      [7:0] n425;
wire      [7:0] n426;
wire      [7:0] n427;
wire      [7:0] n428;
wire      [7:0] n429;
wire      [7:0] n430;
wire      [7:0] n431;
wire      [7:0] n432;
wire      [7:0] n433;
wire      [7:0] n434;
wire      [7:0] n435;
wire      [7:0] n436;
wire      [7:0] n437;
wire      [7:0] n438;
wire      [7:0] n439;
wire      [7:0] n440;
wire      [7:0] n441;
wire      [7:0] n442;
wire      [7:0] n443;
wire      [7:0] n444;
wire      [7:0] n445;
wire      [7:0] n446;
wire      [7:0] n447;
wire      [7:0] n448;
wire      [7:0] n449;
wire      [7:0] n450;
wire      [7:0] n451;
wire      [7:0] n452;
wire      [7:0] n453;
wire      [7:0] n454;
wire      [7:0] n455;
wire      [7:0] n456;
wire      [7:0] n457;
wire      [7:0] n458;
wire     [15:0] n459;
wire     [23:0] n460;
wire     [31:0] n461;
wire     [39:0] n462;
wire     [47:0] n463;
wire     [55:0] n464;
wire     [63:0] n465;
wire     [71:0] n466;
wire     [71:0] n467;
wire     [71:0] n468;
wire     [71:0] n469;
wire     [71:0] n470;
wire     [71:0] n471;
wire     [71:0] n472;
wire     [71:0] n473;
wire     [71:0] n474;
wire     [71:0] n475;
wire     [71:0] n476;
wire     [71:0] n477;
wire     [71:0] n478;
wire     [71:0] n479;
wire     [71:0] n480;
wire     [71:0] n481;
wire     [71:0] n482;
wire            n483;
wire            n484;
wire            n485;
wire            n486;
wire            n487;
wire            n488;
wire            n489;
wire            n490;
wire            n491;
wire            n492;
wire            n493;
wire            n494;
wire            n495;
wire            n496;
wire            n497;
wire            n498;
wire            n499;
wire            n500;
wire            n501;
wire            n502;
wire            n503;
wire            n504;
wire      [7:0] n505;
wire      [7:0] n506;
wire      [7:0] n507;
wire      [7:0] n508;
wire      [7:0] n509;
wire      [7:0] n510;
wire      [7:0] n511;
wire      [7:0] n512;
wire      [7:0] n513;
wire     [15:0] n514;
wire     [23:0] n515;
wire     [31:0] n516;
wire     [39:0] n517;
wire     [47:0] n518;
wire     [55:0] n519;
wire     [63:0] n520;
wire     [71:0] n521;
wire      [7:0] n522;
wire      [7:0] n523;
wire      [7:0] n524;
wire      [7:0] n525;
wire      [7:0] n526;
wire      [7:0] n527;
wire      [7:0] n528;
wire      [7:0] n529;
wire      [7:0] n530;
wire     [15:0] n531;
wire     [23:0] n532;
wire     [31:0] n533;
wire     [39:0] n534;
wire     [47:0] n535;
wire     [55:0] n536;
wire     [63:0] n537;
wire     [71:0] n538;
wire      [7:0] n539;
wire      [7:0] n540;
wire      [7:0] n541;
wire      [7:0] n542;
wire      [7:0] n543;
wire      [7:0] n544;
wire      [7:0] n545;
wire      [7:0] n546;
wire      [7:0] n547;
wire     [15:0] n548;
wire     [23:0] n549;
wire     [31:0] n550;
wire     [39:0] n551;
wire     [47:0] n552;
wire     [55:0] n553;
wire     [63:0] n554;
wire     [71:0] n555;
wire      [7:0] n556;
wire      [7:0] n557;
wire      [7:0] n558;
wire      [7:0] n559;
wire      [7:0] n560;
wire      [7:0] n561;
wire      [7:0] n562;
wire      [7:0] n563;
wire      [7:0] n564;
wire     [15:0] n565;
wire     [23:0] n566;
wire     [31:0] n567;
wire     [39:0] n568;
wire     [47:0] n569;
wire     [55:0] n570;
wire     [63:0] n571;
wire     [71:0] n572;
wire      [7:0] n573;
wire      [7:0] n574;
wire      [7:0] n575;
wire      [7:0] n576;
wire      [7:0] n577;
wire      [7:0] n578;
wire      [7:0] n579;
wire      [7:0] n580;
wire      [7:0] n581;
wire     [15:0] n582;
wire     [23:0] n583;
wire     [31:0] n584;
wire     [39:0] n585;
wire     [47:0] n586;
wire     [55:0] n587;
wire     [63:0] n588;
wire     [71:0] n589;
wire      [7:0] n590;
wire      [7:0] n591;
wire      [7:0] n592;
wire      [7:0] n593;
wire      [7:0] n594;
wire      [7:0] n595;
wire      [7:0] n596;
wire      [7:0] n597;
wire      [7:0] n598;
wire     [15:0] n599;
wire     [23:0] n600;
wire     [31:0] n601;
wire     [39:0] n602;
wire     [47:0] n603;
wire     [55:0] n604;
wire     [63:0] n605;
wire     [71:0] n606;
wire      [7:0] n607;
wire      [7:0] n608;
wire      [7:0] n609;
wire      [7:0] n610;
wire      [7:0] n611;
wire      [7:0] n612;
wire      [7:0] n613;
wire      [7:0] n614;
wire      [7:0] n615;
wire     [15:0] n616;
wire     [23:0] n617;
wire     [31:0] n618;
wire     [39:0] n619;
wire     [47:0] n620;
wire     [55:0] n621;
wire     [63:0] n622;
wire     [71:0] n623;
wire      [7:0] n624;
wire      [7:0] n625;
wire      [7:0] n626;
wire      [7:0] n627;
wire      [7:0] n628;
wire      [7:0] n629;
wire      [7:0] n630;
wire      [7:0] n631;
wire      [7:0] n632;
wire     [15:0] n633;
wire     [23:0] n634;
wire     [31:0] n635;
wire     [39:0] n636;
wire     [47:0] n637;
wire     [55:0] n638;
wire     [63:0] n639;
wire     [71:0] n640;
wire      [7:0] n641;
wire      [7:0] n642;
wire      [7:0] n643;
wire      [7:0] n644;
wire      [7:0] n645;
wire      [7:0] n646;
wire      [7:0] n647;
wire      [7:0] n648;
wire      [7:0] n649;
wire     [15:0] n650;
wire     [23:0] n651;
wire     [31:0] n652;
wire     [39:0] n653;
wire     [47:0] n654;
wire     [55:0] n655;
wire     [63:0] n656;
wire     [71:0] n657;
wire    [143:0] n658;
wire    [215:0] n659;
wire    [287:0] n660;
wire    [359:0] n661;
wire    [431:0] n662;
wire    [503:0] n663;
wire    [575:0] n664;
wire    [647:0] n665;
wire    [647:0] n666;
wire    [647:0] n667;
wire    [647:0] n668;
wire    [647:0] n669;
wire    [647:0] n670;
wire    [647:0] n671;
wire    [647:0] n672;
wire    [647:0] n673;
wire            n674;
wire    [647:0] n675;
wire    [647:0] n676;
wire    [647:0] n677;
wire    [647:0] n678;
wire    [647:0] n679;
wire    [647:0] n680;
wire    [647:0] n681;
wire            n682;
wire            n683;
wire            n684;
wire            n685;
wire            n686;
wire            n687;
wire            n688;
wire            n689;
wire            n690;
wire            n691;
wire            n692;
wire            n693;
wire            n694;
wire            n695;
wire            n696;
wire            n697;
wire            n698;
wire            n699;
wire            n700;
wire            n701;
wire            n702;
wire      [8:0] LB2D_proc_0_addr0;
wire      [7:0] LB2D_proc_0_data0;
wire            n703;
wire            n704;
wire            n705;
wire            n706;
wire            n707;
wire            n708;
wire            n709;
wire            n710;
wire            n711;
wire            n712;
wire            n713;
wire            n714;
wire            n715;
wire            n716;
wire            n717;
wire            n718;
wire            n719;
wire            n720;
wire            n721;
wire            n722;
wire            n723;
wire            n724;
wire      [8:0] LB2D_proc_1_addr0;
wire      [7:0] LB2D_proc_1_data0;
wire            n725;
wire            n726;
wire            n727;
wire      [8:0] LB2D_proc_2_addr0;
wire      [7:0] LB2D_proc_2_data0;
wire            n728;
wire            n729;
wire            n730;
wire      [8:0] LB2D_proc_3_addr0;
wire      [7:0] LB2D_proc_3_data0;
wire            n731;
wire            n732;
wire            n733;
wire      [8:0] LB2D_proc_4_addr0;
wire      [7:0] LB2D_proc_4_data0;
wire            n734;
wire            n735;
wire            n736;
wire      [8:0] LB2D_proc_5_addr0;
wire      [7:0] LB2D_proc_5_data0;
wire            n737;
wire            n738;
wire            n739;
wire      [8:0] LB2D_proc_6_addr0;
wire      [7:0] LB2D_proc_6_data0;
wire            n740;
wire            n741;
wire            n742;
wire      [8:0] LB2D_proc_7_addr0;
wire      [7:0] LB2D_proc_7_data0;
wire            n743;
wire            n744;
wire            n745;
reg      [7:0] LB2D_proc_0[511:0];
reg      [7:0] LB2D_proc_1[511:0];
reg      [7:0] LB2D_proc_2[511:0];
reg      [7:0] LB2D_proc_3[511:0];
reg      [7:0] LB2D_proc_4[511:0];
reg      [7:0] LB2D_proc_5[511:0];
reg      [7:0] LB2D_proc_6[511:0];
reg      [7:0] LB2D_proc_7[511:0];
wire clk;
wire rst;
wire step;
assign n0 =  ( arg_1_TREADY ) == ( 1'd1 )  ;
assign n1 =  ( in_stream_full ) == ( 1'd0 )  ;
assign n2 =  ( n0 ) & ( n1 )  ;
assign n3 =  ( LB1D_it_1 ) == ( 1'd1 )  ;
assign n4 =  ( n2 ) & ( n3 )  ;
assign n5 =  ( LB1D_p_cnt ) == ( 19'd316224 )  ;
assign n6 =  ( n4 ) & ( n5 )  ;
assign n7 =  ( arg_0_TREADY ) == ( 1'd1 )  ;
assign n8 =  ( arg_0_TVALID ) == ( 1'd1 )  ;
assign n9 =  ( n7 ) & ( n8 )  ;
assign n10 =  ( arg_1_TVALID ) == ( 1'd0 )  ;
assign n11 =  ( n9 ) & ( n10 )  ;
assign n12 =  ( arg_1_TVALID ) == ( 1'd1 )  ;
assign n13 =  ( n0 ) & ( n12 )  ;
assign n14 =  ( arg_0_TREADY ) == ( 1'd0 )  ;
assign n15 =  ( n13 ) & ( n14 )  ;
assign n16 =  ( arg_0_TVALID ) == ( 1'd0 )  ;
assign n17 =  ( gb_exit_it_1 ) == ( 1'd0 )  ;
assign n18 =  ( stencil_stream_empty ) == ( 1'd0 )  ;
assign n19 =  ( n17 ) & ( n18 )  ;
assign n20 =  ( gb_exit_it_1 ) == ( 1'd1 )  ;
assign n21 =  ( gb_exit_it_8 ) == ( 1'd0 )  ;
assign n22 =  ( n20 ) & ( n21 )  ;
assign n23 =  ( n19 ) | ( n22 )  ;
assign n24 =  ( n16 ) & ( n23 )  ;
assign n25 =  ( slice_stream_empty ) == ( 1'd0 )  ;
assign n26 =  ( LB2D_shift_x ) != ( 9'd488 )  ;
assign n27 =  ( n25 ) & ( n26 )  ;
assign n28 =  ( stencil_stream_full ) == ( 1'd0 )  ;
assign n29 =  ( LB2D_shift_x ) < ( 9'd8 )  ;
assign n30 =  ( LB2D_shift_x ) > ( 9'd0 )  ;
assign n31 =  ( n29 ) & ( n30 )  ;
assign n32 =  ( n28 ) | ( n31 )  ;
assign n33 =  ( n27 ) & ( n32 )  ;
assign n34 =  ( in_stream_empty ) == ( 1'd0 )  ;
assign n35 =  ( slice_stream_full ) == ( 1'd0 )  ;
assign n36 =  ( LB2D_proc_y ) < ( 10'd8 )  ;
assign n37 =  ( n35 ) | ( n36 )  ;
assign n38 =  ( n34 ) & ( n37 )  ;
assign n39 =  ( arg_1_TREADY ) == ( 1'd0 )  ;
assign n40 =  ( n39 ) & ( n1 )  ;
assign n41 =  ( LB1D_it_1 ) == ( 1'd0 )  ;
assign n42 =  ( n40 ) & ( n41 )  ;
assign n43 =  ( n40 ) & ( n3 )  ;
assign n44 =  ( n43 ) ? ( LB1D_uIn ) : ( LB1D_buff ) ;
assign n45 =  ( n42 ) ? ( LB1D_uIn ) : ( n44 ) ;
assign n46 =  ( n38 ) ? ( LB1D_buff ) : ( n45 ) ;
assign n47 =  ( n33 ) ? ( LB1D_buff ) : ( n46 ) ;
assign n48 =  ( n24 ) ? ( LB1D_buff ) : ( n47 ) ;
assign n49 =  ( n15 ) ? ( LB1D_buff ) : ( n48 ) ;
assign n50 =  ( n11 ) ? ( LB1D_buff ) : ( n49 ) ;
assign n51 =  ( n6 ) ? ( LB1D_uIn ) : ( n50 ) ;
assign n52 =  ( n43 ) ? ( LB1D_in ) : ( LB1D_in ) ;
assign n53 =  ( n42 ) ? ( LB1D_in ) : ( n52 ) ;
assign n54 =  ( n38 ) ? ( LB1D_in ) : ( n53 ) ;
assign n55 =  ( n33 ) ? ( LB1D_in ) : ( n54 ) ;
assign n56 =  ( n24 ) ? ( LB1D_in ) : ( n55 ) ;
assign n57 =  ( n15 ) ? ( arg_1_TDATA ) : ( n56 ) ;
assign n58 =  ( n11 ) ? ( LB1D_in ) : ( n57 ) ;
assign n59 =  ( n6 ) ? ( LB1D_in ) : ( n58 ) ;
assign n60 =  ( n43 ) ? ( 1'd1 ) : ( LB1D_it_1 ) ;
assign n61 =  ( n42 ) ? ( 1'd1 ) : ( n60 ) ;
assign n62 =  ( n6 ) ? ( 1'd0 ) : ( n61 ) ;
assign n63 =  ( LB1D_p_cnt ) + ( 19'd1 )  ;
assign n64 =  ( n43 ) ? ( n63 ) : ( LB1D_p_cnt ) ;
assign n65 =  ( n42 ) ? ( n63 ) : ( n64 ) ;
assign n66 =  ( n38 ) ? ( LB1D_p_cnt ) : ( n65 ) ;
assign n67 =  ( n33 ) ? ( LB1D_p_cnt ) : ( n66 ) ;
assign n68 =  ( n24 ) ? ( LB1D_p_cnt ) : ( n67 ) ;
assign n69 =  ( n15 ) ? ( LB1D_p_cnt ) : ( n68 ) ;
assign n70 =  ( n11 ) ? ( LB1D_p_cnt ) : ( n69 ) ;
assign n71 =  ( n6 ) ? ( 19'd0 ) : ( n70 ) ;
assign n72 =  ( n43 ) ? ( LB1D_in ) : ( LB1D_uIn ) ;
assign n73 =  ( n42 ) ? ( LB1D_in ) : ( n72 ) ;
assign n74 =  ( n38 ) ? ( LB1D_uIn ) : ( n73 ) ;
assign n75 =  ( n33 ) ? ( LB1D_uIn ) : ( n74 ) ;
assign n76 =  ( n24 ) ? ( LB1D_uIn ) : ( n75 ) ;
assign n77 =  ( n15 ) ? ( LB1D_uIn ) : ( n76 ) ;
assign n78 =  ( n6 ) ? ( LB1D_in ) : ( n77 ) ;
assign n79 =  ( LB2D_proc_x ) == ( 9'd488 )  ;
assign n80 =  ( LB2D_proc_w ) == ( 64'd7 )  ;
assign n81 =  ( LB2D_proc_w ) + ( 64'd1 )  ;
assign n82 =  ( n80 ) ? ( 64'd0 ) : ( n81 ) ;
assign n83 =  ( n79 ) ? ( n82 ) : ( LB2D_proc_w ) ;
assign n84 =  ( n43 ) ? ( LB2D_proc_w ) : ( LB2D_proc_w ) ;
assign n85 =  ( n38 ) ? ( n83 ) : ( n84 ) ;
assign n86 =  ( n33 ) ? ( LB2D_proc_w ) : ( n85 ) ;
assign n87 =  ( n24 ) ? ( LB2D_proc_w ) : ( n86 ) ;
assign n88 =  ( n15 ) ? ( LB2D_proc_w ) : ( n87 ) ;
assign n89 =  ( n11 ) ? ( LB2D_proc_w ) : ( n88 ) ;
assign n90 =  ( n6 ) ? ( LB2D_proc_w ) : ( n89 ) ;
assign n91 =  ( LB2D_proc_x ) + ( 9'd1 )  ;
assign n92 =  ( n79 ) ? ( 9'd1 ) : ( n91 ) ;
assign n93 =  ( n43 ) ? ( LB2D_proc_x ) : ( LB2D_proc_x ) ;
assign n94 =  ( n38 ) ? ( n92 ) : ( n93 ) ;
assign n95 =  ( n33 ) ? ( LB2D_proc_x ) : ( n94 ) ;
assign n96 =  ( n24 ) ? ( LB2D_proc_x ) : ( n95 ) ;
assign n97 =  ( n15 ) ? ( LB2D_proc_x ) : ( n96 ) ;
assign n98 =  ( n11 ) ? ( LB2D_proc_x ) : ( n97 ) ;
assign n99 =  ( n6 ) ? ( LB2D_proc_x ) : ( n98 ) ;
assign n100 =  ( LB2D_proc_y ) == ( 10'd648 )  ;
assign n101 =  ( LB2D_proc_y ) + ( 10'd1 )  ;
assign n102 =  ( n100 ) ? ( 10'd0 ) : ( n101 ) ;
assign n103 =  ( n79 ) ? ( n102 ) : ( LB2D_proc_y ) ;
assign n104 =  ( n43 ) ? ( LB2D_proc_y ) : ( LB2D_proc_y ) ;
assign n105 =  ( n38 ) ? ( n103 ) : ( n104 ) ;
assign n106 =  ( n33 ) ? ( LB2D_proc_y ) : ( n105 ) ;
assign n107 =  ( n24 ) ? ( LB2D_proc_y ) : ( n106 ) ;
assign n108 =  ( n15 ) ? ( LB2D_proc_y ) : ( n107 ) ;
assign n109 =  ( n11 ) ? ( LB2D_proc_y ) : ( n108 ) ;
assign n110 =  ( n6 ) ? ( LB2D_proc_y ) : ( n109 ) ;
assign n111 =  ( n43 ) ? ( LB2D_shift_0 ) : ( LB2D_shift_0 ) ;
assign n112 =  ( n38 ) ? ( LB2D_shift_0 ) : ( n111 ) ;
assign n113 =  ( n33 ) ? ( LB2D_shift_1 ) : ( n112 ) ;
assign n114 =  ( n24 ) ? ( LB2D_shift_0 ) : ( n113 ) ;
assign n115 =  ( n15 ) ? ( LB2D_shift_0 ) : ( n114 ) ;
assign n116 =  ( n11 ) ? ( LB2D_shift_0 ) : ( n115 ) ;
assign n117 =  ( n6 ) ? ( LB2D_shift_0 ) : ( n116 ) ;
assign n118 =  ( n43 ) ? ( LB2D_shift_1 ) : ( LB2D_shift_1 ) ;
assign n119 =  ( n38 ) ? ( LB2D_shift_1 ) : ( n118 ) ;
assign n120 =  ( n33 ) ? ( LB2D_shift_2 ) : ( n119 ) ;
assign n121 =  ( n24 ) ? ( LB2D_shift_1 ) : ( n120 ) ;
assign n122 =  ( n15 ) ? ( LB2D_shift_1 ) : ( n121 ) ;
assign n123 =  ( n11 ) ? ( LB2D_shift_1 ) : ( n122 ) ;
assign n124 =  ( n6 ) ? ( LB2D_shift_1 ) : ( n123 ) ;
assign n125 =  ( n43 ) ? ( LB2D_shift_2 ) : ( LB2D_shift_2 ) ;
assign n126 =  ( n38 ) ? ( LB2D_shift_2 ) : ( n125 ) ;
assign n127 =  ( n33 ) ? ( LB2D_shift_3 ) : ( n126 ) ;
assign n128 =  ( n24 ) ? ( LB2D_shift_2 ) : ( n127 ) ;
assign n129 =  ( n15 ) ? ( LB2D_shift_2 ) : ( n128 ) ;
assign n130 =  ( n11 ) ? ( LB2D_shift_2 ) : ( n129 ) ;
assign n131 =  ( n6 ) ? ( LB2D_shift_2 ) : ( n130 ) ;
assign n132 =  ( n43 ) ? ( LB2D_shift_3 ) : ( LB2D_shift_3 ) ;
assign n133 =  ( n38 ) ? ( LB2D_shift_3 ) : ( n132 ) ;
assign n134 =  ( n33 ) ? ( LB2D_shift_4 ) : ( n133 ) ;
assign n135 =  ( n24 ) ? ( LB2D_shift_3 ) : ( n134 ) ;
assign n136 =  ( n15 ) ? ( LB2D_shift_3 ) : ( n135 ) ;
assign n137 =  ( n11 ) ? ( LB2D_shift_3 ) : ( n136 ) ;
assign n138 =  ( n6 ) ? ( LB2D_shift_3 ) : ( n137 ) ;
assign n139 =  ( n43 ) ? ( LB2D_shift_4 ) : ( LB2D_shift_4 ) ;
assign n140 =  ( n38 ) ? ( LB2D_shift_4 ) : ( n139 ) ;
assign n141 =  ( n33 ) ? ( LB2D_shift_5 ) : ( n140 ) ;
assign n142 =  ( n24 ) ? ( LB2D_shift_4 ) : ( n141 ) ;
assign n143 =  ( n15 ) ? ( LB2D_shift_4 ) : ( n142 ) ;
assign n144 =  ( n11 ) ? ( LB2D_shift_4 ) : ( n143 ) ;
assign n145 =  ( n6 ) ? ( LB2D_shift_4 ) : ( n144 ) ;
assign n146 =  ( n43 ) ? ( LB2D_shift_5 ) : ( LB2D_shift_5 ) ;
assign n147 =  ( n38 ) ? ( LB2D_shift_5 ) : ( n146 ) ;
assign n148 =  ( n33 ) ? ( LB2D_shift_6 ) : ( n147 ) ;
assign n149 =  ( n24 ) ? ( LB2D_shift_5 ) : ( n148 ) ;
assign n150 =  ( n15 ) ? ( LB2D_shift_5 ) : ( n149 ) ;
assign n151 =  ( n11 ) ? ( LB2D_shift_5 ) : ( n150 ) ;
assign n152 =  ( n6 ) ? ( LB2D_shift_5 ) : ( n151 ) ;
assign n153 =  ( n43 ) ? ( LB2D_shift_6 ) : ( LB2D_shift_6 ) ;
assign n154 =  ( n38 ) ? ( LB2D_shift_6 ) : ( n153 ) ;
assign n155 =  ( n33 ) ? ( LB2D_shift_7 ) : ( n154 ) ;
assign n156 =  ( n24 ) ? ( LB2D_shift_6 ) : ( n155 ) ;
assign n157 =  ( n15 ) ? ( LB2D_shift_6 ) : ( n156 ) ;
assign n158 =  ( n11 ) ? ( LB2D_shift_6 ) : ( n157 ) ;
assign n159 =  ( n6 ) ? ( LB2D_shift_6 ) : ( n158 ) ;
assign n160 =  ( slice_stream_full ) == ( 1'd1 )  ;
assign n161 =  ( n160 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n162 =  ( n43 ) ? ( LB2D_shift_7 ) : ( LB2D_shift_7 ) ;
assign n163 =  ( n38 ) ? ( LB2D_shift_7 ) : ( n162 ) ;
assign n164 =  ( n33 ) ? ( n161 ) : ( n163 ) ;
assign n165 =  ( n24 ) ? ( LB2D_shift_7 ) : ( n164 ) ;
assign n166 =  ( n15 ) ? ( LB2D_shift_7 ) : ( n165 ) ;
assign n167 =  ( n11 ) ? ( LB2D_shift_7 ) : ( n166 ) ;
assign n168 =  ( n6 ) ? ( LB2D_shift_7 ) : ( n167 ) ;
assign n169 =  ( LB2D_shift_x ) == ( 9'd488 )  ;
assign n170 =  ( n25 ) & ( n169 )  ;
assign n171 =  ( n28 ) | ( n29 )  ;
assign n172 =  ( n170 ) & ( n171 )  ;
assign n173 =  ( LB2D_shift_x ) + ( 9'd1 )  ;
assign n174 =  ( n43 ) ? ( LB2D_shift_x ) : ( LB2D_shift_x ) ;
assign n175 =  ( n38 ) ? ( LB2D_shift_x ) : ( n174 ) ;
assign n176 =  ( n33 ) ? ( n173 ) : ( n175 ) ;
assign n177 =  ( n172 ) ? ( 9'd0 ) : ( n176 ) ;
assign n178 =  ( n24 ) ? ( LB2D_shift_x ) : ( n177 ) ;
assign n179 =  ( n15 ) ? ( LB2D_shift_x ) : ( n178 ) ;
assign n180 =  ( n11 ) ? ( LB2D_shift_x ) : ( n179 ) ;
assign n181 =  ( n6 ) ? ( LB2D_shift_x ) : ( n180 ) ;
assign n182 =  ( LB2D_shift_y ) < ( 10'd640 )  ;
assign n183 =  ( LB2D_shift_x ) < ( 9'd488 )  ;
assign n184 =  ( LB2D_shift_y ) + ( 10'd1 )  ;
assign n185 =  ( n183 ) ? ( LB2D_shift_y ) : ( n184 ) ;
assign n186 =  ( n182 ) ? ( n185 ) : ( 10'd640 ) ;
assign n187 =  ( n43 ) ? ( LB2D_shift_y ) : ( LB2D_shift_y ) ;
assign n188 =  ( n38 ) ? ( LB2D_shift_y ) : ( n187 ) ;
assign n189 =  ( n33 ) ? ( n186 ) : ( n188 ) ;
assign n190 =  ( n24 ) ? ( LB2D_shift_y ) : ( n189 ) ;
assign n191 =  ( n15 ) ? ( LB2D_shift_y ) : ( n190 ) ;
assign n192 =  ( n11 ) ? ( LB2D_shift_y ) : ( n191 ) ;
assign n193 =  ( n6 ) ? ( LB2D_shift_y ) : ( n192 ) ;
assign n194 =  ( stencil_stream_full ) == ( 1'd1 )  ;
assign n195 =  ( n194 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_0 ) ;
assign n196 = gb_fun(n195) ;
assign n197 =  ( n43 ) ? ( arg_0_TDATA ) : ( arg_0_TDATA ) ;
assign n198 =  ( n38 ) ? ( arg_0_TDATA ) : ( n197 ) ;
assign n199 =  ( n33 ) ? ( arg_0_TDATA ) : ( n198 ) ;
assign n200 =  ( n24 ) ? ( n196 ) : ( n199 ) ;
assign n201 =  ( n15 ) ? ( arg_0_TDATA ) : ( n200 ) ;
assign n202 =  ( n11 ) ? ( arg_0_TDATA ) : ( n201 ) ;
assign n203 =  ( n6 ) ? ( arg_0_TDATA ) : ( n202 ) ;
assign n204 =  ( gb_pp_it_8 ) == ( 1'd1 )  ;
assign n205 =  ( gb_exit_it_7 ) == ( 1'd0 )  ;
assign n206 =  ( n204 ) & ( n205 )  ;
assign n207 =  ( n206 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n208 =  ( n43 ) ? ( arg_0_TVALID ) : ( arg_0_TVALID ) ;
assign n209 =  ( n38 ) ? ( arg_0_TVALID ) : ( n208 ) ;
assign n210 =  ( n33 ) ? ( arg_0_TVALID ) : ( n209 ) ;
assign n211 =  ( n24 ) ? ( n207 ) : ( n210 ) ;
assign n212 =  ( n15 ) ? ( arg_0_TVALID ) : ( n211 ) ;
assign n213 =  ( n11 ) ? ( 1'd0 ) : ( n212 ) ;
assign n214 =  ( n6 ) ? ( arg_0_TVALID ) : ( n213 ) ;
assign n215 =  ( n43 ) ? ( 1'd1 ) : ( arg_1_TREADY ) ;
assign n216 =  ( n42 ) ? ( 1'd1 ) : ( n215 ) ;
assign n217 =  ( n38 ) ? ( arg_1_TREADY ) : ( n216 ) ;
assign n218 =  ( n33 ) ? ( arg_1_TREADY ) : ( n217 ) ;
assign n219 =  ( n24 ) ? ( arg_1_TREADY ) : ( n218 ) ;
assign n220 =  ( n15 ) ? ( 1'd0 ) : ( n219 ) ;
assign n221 =  ( n11 ) ? ( arg_1_TREADY ) : ( n220 ) ;
assign n222 =  ( n6 ) ? ( 1'd1 ) : ( n221 ) ;
assign n223 =  ( gb_p_cnt ) == ( 19'd307200 )  ;
assign n224 =  ( n223 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n225 =  ( n43 ) ? ( gb_exit_it_1 ) : ( gb_exit_it_1 ) ;
assign n226 =  ( n38 ) ? ( gb_exit_it_1 ) : ( n225 ) ;
assign n227 =  ( n33 ) ? ( gb_exit_it_1 ) : ( n226 ) ;
assign n228 =  ( n24 ) ? ( n224 ) : ( n227 ) ;
assign n229 =  ( n15 ) ? ( gb_exit_it_1 ) : ( n228 ) ;
assign n230 =  ( n11 ) ? ( gb_exit_it_1 ) : ( n229 ) ;
assign n231 =  ( n6 ) ? ( gb_exit_it_1 ) : ( n230 ) ;
assign n232 =  ( n43 ) ? ( gb_exit_it_2 ) : ( gb_exit_it_2 ) ;
assign n233 =  ( n38 ) ? ( gb_exit_it_2 ) : ( n232 ) ;
assign n234 =  ( n33 ) ? ( gb_exit_it_2 ) : ( n233 ) ;
assign n235 =  ( n24 ) ? ( gb_exit_it_1 ) : ( n234 ) ;
assign n236 =  ( n15 ) ? ( gb_exit_it_2 ) : ( n235 ) ;
assign n237 =  ( n11 ) ? ( gb_exit_it_2 ) : ( n236 ) ;
assign n238 =  ( n6 ) ? ( gb_exit_it_2 ) : ( n237 ) ;
assign n239 =  ( n43 ) ? ( gb_exit_it_3 ) : ( gb_exit_it_3 ) ;
assign n240 =  ( n38 ) ? ( gb_exit_it_3 ) : ( n239 ) ;
assign n241 =  ( n33 ) ? ( gb_exit_it_3 ) : ( n240 ) ;
assign n242 =  ( n24 ) ? ( gb_exit_it_2 ) : ( n241 ) ;
assign n243 =  ( n15 ) ? ( gb_exit_it_3 ) : ( n242 ) ;
assign n244 =  ( n11 ) ? ( gb_exit_it_3 ) : ( n243 ) ;
assign n245 =  ( n6 ) ? ( gb_exit_it_3 ) : ( n244 ) ;
assign n246 =  ( n43 ) ? ( gb_exit_it_4 ) : ( gb_exit_it_4 ) ;
assign n247 =  ( n38 ) ? ( gb_exit_it_4 ) : ( n246 ) ;
assign n248 =  ( n33 ) ? ( gb_exit_it_4 ) : ( n247 ) ;
assign n249 =  ( n24 ) ? ( gb_exit_it_3 ) : ( n248 ) ;
assign n250 =  ( n15 ) ? ( gb_exit_it_4 ) : ( n249 ) ;
assign n251 =  ( n11 ) ? ( gb_exit_it_4 ) : ( n250 ) ;
assign n252 =  ( n6 ) ? ( gb_exit_it_4 ) : ( n251 ) ;
assign n253 =  ( n43 ) ? ( gb_exit_it_5 ) : ( gb_exit_it_5 ) ;
assign n254 =  ( n38 ) ? ( gb_exit_it_5 ) : ( n253 ) ;
assign n255 =  ( n33 ) ? ( gb_exit_it_5 ) : ( n254 ) ;
assign n256 =  ( n24 ) ? ( gb_exit_it_4 ) : ( n255 ) ;
assign n257 =  ( n15 ) ? ( gb_exit_it_5 ) : ( n256 ) ;
assign n258 =  ( n11 ) ? ( gb_exit_it_5 ) : ( n257 ) ;
assign n259 =  ( n6 ) ? ( gb_exit_it_5 ) : ( n258 ) ;
assign n260 =  ( n43 ) ? ( gb_exit_it_6 ) : ( gb_exit_it_6 ) ;
assign n261 =  ( n38 ) ? ( gb_exit_it_6 ) : ( n260 ) ;
assign n262 =  ( n33 ) ? ( gb_exit_it_6 ) : ( n261 ) ;
assign n263 =  ( n24 ) ? ( gb_exit_it_5 ) : ( n262 ) ;
assign n264 =  ( n15 ) ? ( gb_exit_it_6 ) : ( n263 ) ;
assign n265 =  ( n11 ) ? ( gb_exit_it_6 ) : ( n264 ) ;
assign n266 =  ( n6 ) ? ( gb_exit_it_6 ) : ( n265 ) ;
assign n267 =  ( n43 ) ? ( gb_exit_it_7 ) : ( gb_exit_it_7 ) ;
assign n268 =  ( n38 ) ? ( gb_exit_it_7 ) : ( n267 ) ;
assign n269 =  ( n33 ) ? ( gb_exit_it_7 ) : ( n268 ) ;
assign n270 =  ( n24 ) ? ( gb_exit_it_6 ) : ( n269 ) ;
assign n271 =  ( n15 ) ? ( gb_exit_it_7 ) : ( n270 ) ;
assign n272 =  ( n11 ) ? ( gb_exit_it_7 ) : ( n271 ) ;
assign n273 =  ( n6 ) ? ( gb_exit_it_7 ) : ( n272 ) ;
assign n274 =  ( n43 ) ? ( gb_exit_it_8 ) : ( gb_exit_it_8 ) ;
assign n275 =  ( n38 ) ? ( gb_exit_it_8 ) : ( n274 ) ;
assign n276 =  ( n33 ) ? ( gb_exit_it_8 ) : ( n275 ) ;
assign n277 =  ( n24 ) ? ( gb_exit_it_7 ) : ( n276 ) ;
assign n278 =  ( n15 ) ? ( gb_exit_it_8 ) : ( n277 ) ;
assign n279 =  ( n11 ) ? ( gb_exit_it_8 ) : ( n278 ) ;
assign n280 =  ( n6 ) ? ( gb_exit_it_8 ) : ( n279 ) ;
assign n281 =  ( gb_p_cnt ) < ( 19'd307200 )  ;
assign n282 =  ( gb_p_cnt ) + ( 19'd1 )  ;
assign n283 =  ( n281 ) ? ( n282 ) : ( 19'd307200 ) ;
assign n284 =  ( n43 ) ? ( gb_p_cnt ) : ( gb_p_cnt ) ;
assign n285 =  ( n38 ) ? ( gb_p_cnt ) : ( n284 ) ;
assign n286 =  ( n33 ) ? ( gb_p_cnt ) : ( n285 ) ;
assign n287 =  ( n24 ) ? ( n283 ) : ( n286 ) ;
assign n288 =  ( n15 ) ? ( gb_p_cnt ) : ( n287 ) ;
assign n289 =  ( n11 ) ? ( gb_p_cnt ) : ( n288 ) ;
assign n290 =  ( n6 ) ? ( gb_p_cnt ) : ( n289 ) ;
assign n291 =  ( n43 ) ? ( gb_pp_it_1 ) : ( gb_pp_it_1 ) ;
assign n292 =  ( n38 ) ? ( gb_pp_it_1 ) : ( n291 ) ;
assign n293 =  ( n33 ) ? ( gb_pp_it_1 ) : ( n292 ) ;
assign n294 =  ( n24 ) ? ( 1'd1 ) : ( n293 ) ;
assign n295 =  ( n15 ) ? ( gb_pp_it_1 ) : ( n294 ) ;
assign n296 =  ( n11 ) ? ( gb_pp_it_1 ) : ( n295 ) ;
assign n297 =  ( n6 ) ? ( gb_pp_it_1 ) : ( n296 ) ;
assign n298 =  ( n43 ) ? ( gb_pp_it_2 ) : ( gb_pp_it_2 ) ;
assign n299 =  ( n38 ) ? ( gb_pp_it_2 ) : ( n298 ) ;
assign n300 =  ( n33 ) ? ( gb_pp_it_2 ) : ( n299 ) ;
assign n301 =  ( n24 ) ? ( gb_pp_it_1 ) : ( n300 ) ;
assign n302 =  ( n15 ) ? ( gb_pp_it_2 ) : ( n301 ) ;
assign n303 =  ( n11 ) ? ( gb_pp_it_2 ) : ( n302 ) ;
assign n304 =  ( n6 ) ? ( gb_pp_it_2 ) : ( n303 ) ;
assign n305 =  ( n43 ) ? ( gb_pp_it_3 ) : ( gb_pp_it_3 ) ;
assign n306 =  ( n38 ) ? ( gb_pp_it_3 ) : ( n305 ) ;
assign n307 =  ( n33 ) ? ( gb_pp_it_3 ) : ( n306 ) ;
assign n308 =  ( n24 ) ? ( gb_pp_it_2 ) : ( n307 ) ;
assign n309 =  ( n15 ) ? ( gb_pp_it_3 ) : ( n308 ) ;
assign n310 =  ( n11 ) ? ( gb_pp_it_3 ) : ( n309 ) ;
assign n311 =  ( n6 ) ? ( gb_pp_it_3 ) : ( n310 ) ;
assign n312 =  ( n43 ) ? ( gb_pp_it_4 ) : ( gb_pp_it_4 ) ;
assign n313 =  ( n38 ) ? ( gb_pp_it_4 ) : ( n312 ) ;
assign n314 =  ( n33 ) ? ( gb_pp_it_4 ) : ( n313 ) ;
assign n315 =  ( n24 ) ? ( gb_pp_it_3 ) : ( n314 ) ;
assign n316 =  ( n15 ) ? ( gb_pp_it_4 ) : ( n315 ) ;
assign n317 =  ( n11 ) ? ( gb_pp_it_4 ) : ( n316 ) ;
assign n318 =  ( n6 ) ? ( gb_pp_it_4 ) : ( n317 ) ;
assign n319 =  ( n43 ) ? ( gb_pp_it_5 ) : ( gb_pp_it_5 ) ;
assign n320 =  ( n38 ) ? ( gb_pp_it_5 ) : ( n319 ) ;
assign n321 =  ( n33 ) ? ( gb_pp_it_5 ) : ( n320 ) ;
assign n322 =  ( n24 ) ? ( gb_pp_it_4 ) : ( n321 ) ;
assign n323 =  ( n15 ) ? ( gb_pp_it_5 ) : ( n322 ) ;
assign n324 =  ( n11 ) ? ( gb_pp_it_5 ) : ( n323 ) ;
assign n325 =  ( n6 ) ? ( gb_pp_it_5 ) : ( n324 ) ;
assign n326 =  ( n43 ) ? ( gb_pp_it_6 ) : ( gb_pp_it_6 ) ;
assign n327 =  ( n38 ) ? ( gb_pp_it_6 ) : ( n326 ) ;
assign n328 =  ( n33 ) ? ( gb_pp_it_6 ) : ( n327 ) ;
assign n329 =  ( n24 ) ? ( gb_pp_it_5 ) : ( n328 ) ;
assign n330 =  ( n15 ) ? ( gb_pp_it_6 ) : ( n329 ) ;
assign n331 =  ( n11 ) ? ( gb_pp_it_6 ) : ( n330 ) ;
assign n332 =  ( n6 ) ? ( gb_pp_it_6 ) : ( n331 ) ;
assign n333 =  ( n43 ) ? ( gb_pp_it_7 ) : ( gb_pp_it_7 ) ;
assign n334 =  ( n38 ) ? ( gb_pp_it_7 ) : ( n333 ) ;
assign n335 =  ( n33 ) ? ( gb_pp_it_7 ) : ( n334 ) ;
assign n336 =  ( n24 ) ? ( gb_pp_it_6 ) : ( n335 ) ;
assign n337 =  ( n15 ) ? ( gb_pp_it_7 ) : ( n336 ) ;
assign n338 =  ( n11 ) ? ( gb_pp_it_7 ) : ( n337 ) ;
assign n339 =  ( n6 ) ? ( gb_pp_it_7 ) : ( n338 ) ;
assign n340 =  ( n43 ) ? ( gb_pp_it_8 ) : ( gb_pp_it_8 ) ;
assign n341 =  ( n38 ) ? ( gb_pp_it_8 ) : ( n340 ) ;
assign n342 =  ( n33 ) ? ( gb_pp_it_8 ) : ( n341 ) ;
assign n343 =  ( n24 ) ? ( gb_pp_it_7 ) : ( n342 ) ;
assign n344 =  ( n15 ) ? ( gb_pp_it_8 ) : ( n343 ) ;
assign n345 =  ( n11 ) ? ( gb_pp_it_8 ) : ( n344 ) ;
assign n346 =  ( n6 ) ? ( gb_pp_it_8 ) : ( n345 ) ;
assign n347 =  ( n43 ) ? ( gb_pp_it_9 ) : ( gb_pp_it_9 ) ;
assign n348 =  ( n38 ) ? ( gb_pp_it_9 ) : ( n347 ) ;
assign n349 =  ( n33 ) ? ( gb_pp_it_9 ) : ( n348 ) ;
assign n350 =  ( n24 ) ? ( gb_pp_it_8 ) : ( n349 ) ;
assign n351 =  ( n15 ) ? ( gb_pp_it_9 ) : ( n350 ) ;
assign n352 =  ( n11 ) ? ( gb_pp_it_9 ) : ( n351 ) ;
assign n353 =  ( n6 ) ? ( gb_pp_it_9 ) : ( n352 ) ;
assign n354 =  ( n43 ) ? ( LB1D_uIn ) : ( in_stream_buff_0 ) ;
assign n355 =  ( n38 ) ? ( in_stream_buff_0 ) : ( n354 ) ;
assign n356 =  ( n33 ) ? ( in_stream_buff_0 ) : ( n355 ) ;
assign n357 =  ( n24 ) ? ( in_stream_buff_0 ) : ( n356 ) ;
assign n358 =  ( n15 ) ? ( in_stream_buff_0 ) : ( n357 ) ;
assign n359 =  ( n11 ) ? ( in_stream_buff_0 ) : ( n358 ) ;
assign n360 =  ( n6 ) ? ( LB1D_uIn ) : ( n359 ) ;
assign n361 =  ( n43 ) ? ( in_stream_buff_0 ) : ( in_stream_buff_1 ) ;
assign n362 =  ( n38 ) ? ( in_stream_buff_1 ) : ( n361 ) ;
assign n363 =  ( n33 ) ? ( in_stream_buff_1 ) : ( n362 ) ;
assign n364 =  ( n24 ) ? ( in_stream_buff_1 ) : ( n363 ) ;
assign n365 =  ( n15 ) ? ( in_stream_buff_1 ) : ( n364 ) ;
assign n366 =  ( n11 ) ? ( in_stream_buff_1 ) : ( n365 ) ;
assign n367 =  ( n6 ) ? ( in_stream_buff_0 ) : ( n366 ) ;
assign n368 =  ( in_stream_full ) == ( 1'd1 )  ;
assign n369 =  ( n368 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n370 =  ( n43 ) ? ( 1'd0 ) : ( in_stream_empty ) ;
assign n371 =  ( n38 ) ? ( n369 ) : ( n370 ) ;
assign n372 =  ( n33 ) ? ( in_stream_empty ) : ( n371 ) ;
assign n373 =  ( n24 ) ? ( in_stream_empty ) : ( n372 ) ;
assign n374 =  ( n15 ) ? ( in_stream_empty ) : ( n373 ) ;
assign n375 =  ( n11 ) ? ( in_stream_empty ) : ( n374 ) ;
assign n376 =  ( n6 ) ? ( 1'd0 ) : ( n375 ) ;
assign n377 =  ( in_stream_empty ) == ( 1'd1 )  ;
assign n378 =  ( n377 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n379 =  ( n43 ) ? ( n378 ) : ( in_stream_full ) ;
assign n380 =  ( n38 ) ? ( 1'd0 ) : ( n379 ) ;
assign n381 =  ( n33 ) ? ( in_stream_full ) : ( n380 ) ;
assign n382 =  ( n24 ) ? ( in_stream_full ) : ( n381 ) ;
assign n383 =  ( n15 ) ? ( in_stream_full ) : ( n382 ) ;
assign n384 =  ( n11 ) ? ( in_stream_full ) : ( n383 ) ;
assign n385 =  ( n6 ) ? ( n378 ) : ( n384 ) ;
assign n386 =  ( n368 ) ? ( in_stream_buff_1 ) : ( in_stream_buff_0 ) ;
assign n387 =  ( LB2D_proc_w ) == ( 64'd0 )  ;
assign n388 =  ( LB2D_proc_x ) - ( 9'd1 )  ;
assign n389 =  (  LB2D_proc_7 [ n388 ] )  ;
assign n390 =  ( LB2D_proc_w ) == ( 64'd1 )  ;
assign n391 =  (  LB2D_proc_0 [ n388 ] )  ;
assign n392 =  ( LB2D_proc_w ) == ( 64'd2 )  ;
assign n393 =  (  LB2D_proc_1 [ n388 ] )  ;
assign n394 =  ( LB2D_proc_w ) == ( 64'd3 )  ;
assign n395 =  (  LB2D_proc_2 [ n388 ] )  ;
assign n396 =  ( LB2D_proc_w ) == ( 64'd4 )  ;
assign n397 =  (  LB2D_proc_3 [ n388 ] )  ;
assign n398 =  ( LB2D_proc_w ) == ( 64'd5 )  ;
assign n399 =  (  LB2D_proc_4 [ n388 ] )  ;
assign n400 =  ( LB2D_proc_w ) == ( 64'd6 )  ;
assign n401 =  (  LB2D_proc_5 [ n388 ] )  ;
assign n402 =  (  LB2D_proc_6 [ n388 ] )  ;
assign n403 =  ( n400 ) ? ( n401 ) : ( n402 ) ;
assign n404 =  ( n398 ) ? ( n399 ) : ( n403 ) ;
assign n405 =  ( n396 ) ? ( n397 ) : ( n404 ) ;
assign n406 =  ( n394 ) ? ( n395 ) : ( n405 ) ;
assign n407 =  ( n392 ) ? ( n393 ) : ( n406 ) ;
assign n408 =  ( n390 ) ? ( n391 ) : ( n407 ) ;
assign n409 =  ( n387 ) ? ( n389 ) : ( n408 ) ;
assign n410 =  ( n400 ) ? ( n399 ) : ( n401 ) ;
assign n411 =  ( n398 ) ? ( n397 ) : ( n410 ) ;
assign n412 =  ( n396 ) ? ( n395 ) : ( n411 ) ;
assign n413 =  ( n394 ) ? ( n393 ) : ( n412 ) ;
assign n414 =  ( n392 ) ? ( n391 ) : ( n413 ) ;
assign n415 =  ( n390 ) ? ( n389 ) : ( n414 ) ;
assign n416 =  ( n387 ) ? ( n402 ) : ( n415 ) ;
assign n417 =  ( n400 ) ? ( n397 ) : ( n399 ) ;
assign n418 =  ( n398 ) ? ( n395 ) : ( n417 ) ;
assign n419 =  ( n396 ) ? ( n393 ) : ( n418 ) ;
assign n420 =  ( n394 ) ? ( n391 ) : ( n419 ) ;
assign n421 =  ( n392 ) ? ( n389 ) : ( n420 ) ;
assign n422 =  ( n390 ) ? ( n402 ) : ( n421 ) ;
assign n423 =  ( n387 ) ? ( n401 ) : ( n422 ) ;
assign n424 =  ( n400 ) ? ( n395 ) : ( n397 ) ;
assign n425 =  ( n398 ) ? ( n393 ) : ( n424 ) ;
assign n426 =  ( n396 ) ? ( n391 ) : ( n425 ) ;
assign n427 =  ( n394 ) ? ( n389 ) : ( n426 ) ;
assign n428 =  ( n392 ) ? ( n402 ) : ( n427 ) ;
assign n429 =  ( n390 ) ? ( n401 ) : ( n428 ) ;
assign n430 =  ( n387 ) ? ( n399 ) : ( n429 ) ;
assign n431 =  ( n400 ) ? ( n393 ) : ( n395 ) ;
assign n432 =  ( n398 ) ? ( n391 ) : ( n431 ) ;
assign n433 =  ( n396 ) ? ( n389 ) : ( n432 ) ;
assign n434 =  ( n394 ) ? ( n402 ) : ( n433 ) ;
assign n435 =  ( n392 ) ? ( n401 ) : ( n434 ) ;
assign n436 =  ( n390 ) ? ( n399 ) : ( n435 ) ;
assign n437 =  ( n387 ) ? ( n397 ) : ( n436 ) ;
assign n438 =  ( n400 ) ? ( n391 ) : ( n393 ) ;
assign n439 =  ( n398 ) ? ( n389 ) : ( n438 ) ;
assign n440 =  ( n396 ) ? ( n402 ) : ( n439 ) ;
assign n441 =  ( n394 ) ? ( n401 ) : ( n440 ) ;
assign n442 =  ( n392 ) ? ( n399 ) : ( n441 ) ;
assign n443 =  ( n390 ) ? ( n397 ) : ( n442 ) ;
assign n444 =  ( n387 ) ? ( n395 ) : ( n443 ) ;
assign n445 =  ( n400 ) ? ( n389 ) : ( n391 ) ;
assign n446 =  ( n398 ) ? ( n402 ) : ( n445 ) ;
assign n447 =  ( n396 ) ? ( n401 ) : ( n446 ) ;
assign n448 =  ( n394 ) ? ( n399 ) : ( n447 ) ;
assign n449 =  ( n392 ) ? ( n397 ) : ( n448 ) ;
assign n450 =  ( n390 ) ? ( n395 ) : ( n449 ) ;
assign n451 =  ( n387 ) ? ( n393 ) : ( n450 ) ;
assign n452 =  ( n400 ) ? ( n402 ) : ( n389 ) ;
assign n453 =  ( n398 ) ? ( n401 ) : ( n452 ) ;
assign n454 =  ( n396 ) ? ( n399 ) : ( n453 ) ;
assign n455 =  ( n394 ) ? ( n397 ) : ( n454 ) ;
assign n456 =  ( n392 ) ? ( n395 ) : ( n455 ) ;
assign n457 =  ( n390 ) ? ( n393 ) : ( n456 ) ;
assign n458 =  ( n387 ) ? ( n391 ) : ( n457 ) ;
assign n459 =  { ( n451 ) , ( n458 ) }  ;
assign n460 =  { ( n444 ) , ( n459 ) }  ;
assign n461 =  { ( n437 ) , ( n460 ) }  ;
assign n462 =  { ( n430 ) , ( n461 ) }  ;
assign n463 =  { ( n423 ) , ( n462 ) }  ;
assign n464 =  { ( n416 ) , ( n463 ) }  ;
assign n465 =  { ( n409 ) , ( n464 ) }  ;
assign n466 =  { ( n386 ) , ( n465 ) }  ;
assign n467 =  ( n36 ) ? ( slice_stream_buff_0 ) : ( n466 ) ;
assign n468 =  ( n43 ) ? ( slice_stream_buff_0 ) : ( slice_stream_buff_0 ) ;
assign n469 =  ( n38 ) ? ( n467 ) : ( n468 ) ;
assign n470 =  ( n33 ) ? ( slice_stream_buff_0 ) : ( n469 ) ;
assign n471 =  ( n24 ) ? ( slice_stream_buff_0 ) : ( n470 ) ;
assign n472 =  ( n15 ) ? ( slice_stream_buff_0 ) : ( n471 ) ;
assign n473 =  ( n11 ) ? ( slice_stream_buff_0 ) : ( n472 ) ;
assign n474 =  ( n6 ) ? ( slice_stream_buff_0 ) : ( n473 ) ;
assign n475 =  ( n36 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n476 =  ( n43 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_1 ) ;
assign n477 =  ( n38 ) ? ( n475 ) : ( n476 ) ;
assign n478 =  ( n33 ) ? ( slice_stream_buff_1 ) : ( n477 ) ;
assign n479 =  ( n24 ) ? ( slice_stream_buff_1 ) : ( n478 ) ;
assign n480 =  ( n15 ) ? ( slice_stream_buff_1 ) : ( n479 ) ;
assign n481 =  ( n11 ) ? ( slice_stream_buff_1 ) : ( n480 ) ;
assign n482 =  ( n6 ) ? ( slice_stream_buff_1 ) : ( n481 ) ;
assign n483 =  ( n160 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n484 =  ( n36 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n485 =  ( n43 ) ? ( slice_stream_empty ) : ( slice_stream_empty ) ;
assign n486 =  ( n38 ) ? ( n484 ) : ( n485 ) ;
assign n487 =  ( n33 ) ? ( n483 ) : ( n486 ) ;
assign n488 =  ( n24 ) ? ( slice_stream_empty ) : ( n487 ) ;
assign n489 =  ( n15 ) ? ( slice_stream_empty ) : ( n488 ) ;
assign n490 =  ( n11 ) ? ( slice_stream_empty ) : ( n489 ) ;
assign n491 =  ( n6 ) ? ( slice_stream_empty ) : ( n490 ) ;
assign n492 =  ( slice_stream_empty ) == ( 1'd1 )  ;
assign n493 =  ( n492 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n494 =  ( n36 ) ? ( 1'd0 ) : ( n493 ) ;
assign n495 =  ( n43 ) ? ( slice_stream_full ) : ( slice_stream_full ) ;
assign n496 =  ( n38 ) ? ( n494 ) : ( n495 ) ;
assign n497 =  ( n33 ) ? ( 1'd0 ) : ( n496 ) ;
assign n498 =  ( n24 ) ? ( slice_stream_full ) : ( n497 ) ;
assign n499 =  ( n15 ) ? ( slice_stream_full ) : ( n498 ) ;
assign n500 =  ( n11 ) ? ( slice_stream_full ) : ( n499 ) ;
assign n501 =  ( n6 ) ? ( slice_stream_full ) : ( n500 ) ;
assign n502 =  ( LB2D_shift_x ) >= ( 9'd8 )  ;
assign n503 =  ( LB2D_shift_x ) == ( 9'd0 )  ;
assign n504 =  ( n502 ) | ( n503 )  ;
assign n505 = n161[71:64] ;
assign n506 = LB2D_shift_7[71:64] ;
assign n507 = LB2D_shift_6[71:64] ;
assign n508 = LB2D_shift_5[71:64] ;
assign n509 = LB2D_shift_4[71:64] ;
assign n510 = LB2D_shift_3[71:64] ;
assign n511 = LB2D_shift_2[71:64] ;
assign n512 = LB2D_shift_1[71:64] ;
assign n513 = LB2D_shift_0[71:64] ;
assign n514 =  { ( n512 ) , ( n513 ) }  ;
assign n515 =  { ( n511 ) , ( n514 ) }  ;
assign n516 =  { ( n510 ) , ( n515 ) }  ;
assign n517 =  { ( n509 ) , ( n516 ) }  ;
assign n518 =  { ( n508 ) , ( n517 ) }  ;
assign n519 =  { ( n507 ) , ( n518 ) }  ;
assign n520 =  { ( n506 ) , ( n519 ) }  ;
assign n521 =  { ( n505 ) , ( n520 ) }  ;
assign n522 = n161[63:56] ;
assign n523 = LB2D_shift_7[63:56] ;
assign n524 = LB2D_shift_6[63:56] ;
assign n525 = LB2D_shift_5[63:56] ;
assign n526 = LB2D_shift_4[63:56] ;
assign n527 = LB2D_shift_3[63:56] ;
assign n528 = LB2D_shift_2[63:56] ;
assign n529 = LB2D_shift_1[63:56] ;
assign n530 = LB2D_shift_0[63:56] ;
assign n531 =  { ( n529 ) , ( n530 ) }  ;
assign n532 =  { ( n528 ) , ( n531 ) }  ;
assign n533 =  { ( n527 ) , ( n532 ) }  ;
assign n534 =  { ( n526 ) , ( n533 ) }  ;
assign n535 =  { ( n525 ) , ( n534 ) }  ;
assign n536 =  { ( n524 ) , ( n535 ) }  ;
assign n537 =  { ( n523 ) , ( n536 ) }  ;
assign n538 =  { ( n522 ) , ( n537 ) }  ;
assign n539 = n161[55:48] ;
assign n540 = LB2D_shift_7[55:48] ;
assign n541 = LB2D_shift_6[55:48] ;
assign n542 = LB2D_shift_5[55:48] ;
assign n543 = LB2D_shift_4[55:48] ;
assign n544 = LB2D_shift_3[55:48] ;
assign n545 = LB2D_shift_2[55:48] ;
assign n546 = LB2D_shift_1[55:48] ;
assign n547 = LB2D_shift_0[55:48] ;
assign n548 =  { ( n546 ) , ( n547 ) }  ;
assign n549 =  { ( n545 ) , ( n548 ) }  ;
assign n550 =  { ( n544 ) , ( n549 ) }  ;
assign n551 =  { ( n543 ) , ( n550 ) }  ;
assign n552 =  { ( n542 ) , ( n551 ) }  ;
assign n553 =  { ( n541 ) , ( n552 ) }  ;
assign n554 =  { ( n540 ) , ( n553 ) }  ;
assign n555 =  { ( n539 ) , ( n554 ) }  ;
assign n556 = n161[47:40] ;
assign n557 = LB2D_shift_7[47:40] ;
assign n558 = LB2D_shift_6[47:40] ;
assign n559 = LB2D_shift_5[47:40] ;
assign n560 = LB2D_shift_4[47:40] ;
assign n561 = LB2D_shift_3[47:40] ;
assign n562 = LB2D_shift_2[47:40] ;
assign n563 = LB2D_shift_1[47:40] ;
assign n564 = LB2D_shift_0[47:40] ;
assign n565 =  { ( n563 ) , ( n564 ) }  ;
assign n566 =  { ( n562 ) , ( n565 ) }  ;
assign n567 =  { ( n561 ) , ( n566 ) }  ;
assign n568 =  { ( n560 ) , ( n567 ) }  ;
assign n569 =  { ( n559 ) , ( n568 ) }  ;
assign n570 =  { ( n558 ) , ( n569 ) }  ;
assign n571 =  { ( n557 ) , ( n570 ) }  ;
assign n572 =  { ( n556 ) , ( n571 ) }  ;
assign n573 = n161[39:32] ;
assign n574 = LB2D_shift_7[39:32] ;
assign n575 = LB2D_shift_6[39:32] ;
assign n576 = LB2D_shift_5[39:32] ;
assign n577 = LB2D_shift_4[39:32] ;
assign n578 = LB2D_shift_3[39:32] ;
assign n579 = LB2D_shift_2[39:32] ;
assign n580 = LB2D_shift_1[39:32] ;
assign n581 = LB2D_shift_0[39:32] ;
assign n582 =  { ( n580 ) , ( n581 ) }  ;
assign n583 =  { ( n579 ) , ( n582 ) }  ;
assign n584 =  { ( n578 ) , ( n583 ) }  ;
assign n585 =  { ( n577 ) , ( n584 ) }  ;
assign n586 =  { ( n576 ) , ( n585 ) }  ;
assign n587 =  { ( n575 ) , ( n586 ) }  ;
assign n588 =  { ( n574 ) , ( n587 ) }  ;
assign n589 =  { ( n573 ) , ( n588 ) }  ;
assign n590 = n161[31:24] ;
assign n591 = LB2D_shift_7[31:24] ;
assign n592 = LB2D_shift_6[31:24] ;
assign n593 = LB2D_shift_5[31:24] ;
assign n594 = LB2D_shift_4[31:24] ;
assign n595 = LB2D_shift_3[31:24] ;
assign n596 = LB2D_shift_2[31:24] ;
assign n597 = LB2D_shift_1[31:24] ;
assign n598 = LB2D_shift_0[31:24] ;
assign n599 =  { ( n597 ) , ( n598 ) }  ;
assign n600 =  { ( n596 ) , ( n599 ) }  ;
assign n601 =  { ( n595 ) , ( n600 ) }  ;
assign n602 =  { ( n594 ) , ( n601 ) }  ;
assign n603 =  { ( n593 ) , ( n602 ) }  ;
assign n604 =  { ( n592 ) , ( n603 ) }  ;
assign n605 =  { ( n591 ) , ( n604 ) }  ;
assign n606 =  { ( n590 ) , ( n605 ) }  ;
assign n607 = n161[23:16] ;
assign n608 = LB2D_shift_7[23:16] ;
assign n609 = LB2D_shift_6[23:16] ;
assign n610 = LB2D_shift_5[23:16] ;
assign n611 = LB2D_shift_4[23:16] ;
assign n612 = LB2D_shift_3[23:16] ;
assign n613 = LB2D_shift_2[23:16] ;
assign n614 = LB2D_shift_1[23:16] ;
assign n615 = LB2D_shift_0[23:16] ;
assign n616 =  { ( n614 ) , ( n615 ) }  ;
assign n617 =  { ( n613 ) , ( n616 ) }  ;
assign n618 =  { ( n612 ) , ( n617 ) }  ;
assign n619 =  { ( n611 ) , ( n618 ) }  ;
assign n620 =  { ( n610 ) , ( n619 ) }  ;
assign n621 =  { ( n609 ) , ( n620 ) }  ;
assign n622 =  { ( n608 ) , ( n621 ) }  ;
assign n623 =  { ( n607 ) , ( n622 ) }  ;
assign n624 = n161[15:8] ;
assign n625 = LB2D_shift_7[15:8] ;
assign n626 = LB2D_shift_6[15:8] ;
assign n627 = LB2D_shift_5[15:8] ;
assign n628 = LB2D_shift_4[15:8] ;
assign n629 = LB2D_shift_3[15:8] ;
assign n630 = LB2D_shift_2[15:8] ;
assign n631 = LB2D_shift_1[15:8] ;
assign n632 = LB2D_shift_0[15:8] ;
assign n633 =  { ( n631 ) , ( n632 ) }  ;
assign n634 =  { ( n630 ) , ( n633 ) }  ;
assign n635 =  { ( n629 ) , ( n634 ) }  ;
assign n636 =  { ( n628 ) , ( n635 ) }  ;
assign n637 =  { ( n627 ) , ( n636 ) }  ;
assign n638 =  { ( n626 ) , ( n637 ) }  ;
assign n639 =  { ( n625 ) , ( n638 ) }  ;
assign n640 =  { ( n624 ) , ( n639 ) }  ;
assign n641 = n161[7:0] ;
assign n642 = LB2D_shift_7[7:0] ;
assign n643 = LB2D_shift_6[7:0] ;
assign n644 = LB2D_shift_5[7:0] ;
assign n645 = LB2D_shift_4[7:0] ;
assign n646 = LB2D_shift_3[7:0] ;
assign n647 = LB2D_shift_2[7:0] ;
assign n648 = LB2D_shift_1[7:0] ;
assign n649 = LB2D_shift_0[7:0] ;
assign n650 =  { ( n648 ) , ( n649 ) }  ;
assign n651 =  { ( n647 ) , ( n650 ) }  ;
assign n652 =  { ( n646 ) , ( n651 ) }  ;
assign n653 =  { ( n645 ) , ( n652 ) }  ;
assign n654 =  { ( n644 ) , ( n653 ) }  ;
assign n655 =  { ( n643 ) , ( n654 ) }  ;
assign n656 =  { ( n642 ) , ( n655 ) }  ;
assign n657 =  { ( n641 ) , ( n656 ) }  ;
assign n658 =  { ( n640 ) , ( n657 ) }  ;
assign n659 =  { ( n623 ) , ( n658 ) }  ;
assign n660 =  { ( n606 ) , ( n659 ) }  ;
assign n661 =  { ( n589 ) , ( n660 ) }  ;
assign n662 =  { ( n572 ) , ( n661 ) }  ;
assign n663 =  { ( n555 ) , ( n662 ) }  ;
assign n664 =  { ( n538 ) , ( n663 ) }  ;
assign n665 =  { ( n521 ) , ( n664 ) }  ;
assign n666 =  ( n504 ) ? ( n665 ) : ( stencil_stream_buff_0 ) ;
assign n667 =  ( n43 ) ? ( stencil_stream_buff_0 ) : ( stencil_stream_buff_0 ) ;
assign n668 =  ( n38 ) ? ( stencil_stream_buff_0 ) : ( n667 ) ;
assign n669 =  ( n33 ) ? ( n666 ) : ( n668 ) ;
assign n670 =  ( n24 ) ? ( stencil_stream_buff_0 ) : ( n669 ) ;
assign n671 =  ( n15 ) ? ( stencil_stream_buff_0 ) : ( n670 ) ;
assign n672 =  ( n11 ) ? ( stencil_stream_buff_0 ) : ( n671 ) ;
assign n673 =  ( n6 ) ? ( stencil_stream_buff_0 ) : ( n672 ) ;
assign n674 =  ( n33 ) & ( n504 )  ;
assign n675 =  ( n43 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_1 ) ;
assign n676 =  ( n38 ) ? ( stencil_stream_buff_1 ) : ( n675 ) ;
assign n677 =  ( n674 ) ? ( stencil_stream_buff_0 ) : ( n676 ) ;
assign n678 =  ( n24 ) ? ( stencil_stream_buff_1 ) : ( n677 ) ;
assign n679 =  ( n15 ) ? ( stencil_stream_buff_1 ) : ( n678 ) ;
assign n680 =  ( n11 ) ? ( stencil_stream_buff_1 ) : ( n679 ) ;
assign n681 =  ( n6 ) ? ( stencil_stream_buff_1 ) : ( n680 ) ;
assign n682 =  ( n194 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n683 = ~ ( n504 ) ;
assign n684 =  ( n683 ) ? ( stencil_stream_empty ) : ( 1'd0 ) ;
assign n685 =  ( n43 ) ? ( stencil_stream_empty ) : ( stencil_stream_empty ) ;
assign n686 =  ( n38 ) ? ( stencil_stream_empty ) : ( n685 ) ;
assign n687 =  ( n33 ) ? ( n684 ) : ( n686 ) ;
assign n688 =  ( n24 ) ? ( n682 ) : ( n687 ) ;
assign n689 =  ( n15 ) ? ( stencil_stream_empty ) : ( n688 ) ;
assign n690 =  ( n11 ) ? ( stencil_stream_empty ) : ( n689 ) ;
assign n691 =  ( n6 ) ? ( stencil_stream_empty ) : ( n690 ) ;
assign n692 =  ( n20 ) ? ( 1'd0 ) : ( 1'd0 ) ;
assign n693 =  ( stencil_stream_empty ) == ( 1'd1 )  ;
assign n694 =  ( n693 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n695 =  ( n683 ) ? ( stencil_stream_full ) : ( n694 ) ;
assign n696 =  ( n43 ) ? ( stencil_stream_full ) : ( stencil_stream_full ) ;
assign n697 =  ( n38 ) ? ( stencil_stream_full ) : ( n696 ) ;
assign n698 =  ( n33 ) ? ( n695 ) : ( n697 ) ;
assign n699 =  ( n24 ) ? ( n692 ) : ( n698 ) ;
assign n700 =  ( n15 ) ? ( stencil_stream_full ) : ( n699 ) ;
assign n701 =  ( n11 ) ? ( stencil_stream_full ) : ( n700 ) ;
assign n702 =  ( n6 ) ? ( stencil_stream_full ) : ( n701 ) ;
assign n703 = ~ ( n6 ) ;
assign n704 = ~ ( n11 ) ;
assign n705 =  ( n703 ) & ( n704 )  ;
assign n706 = ~ ( n15 ) ;
assign n707 =  ( n705 ) & ( n706 )  ;
assign n708 = ~ ( n24 ) ;
assign n709 =  ( n707 ) & ( n708 )  ;
assign n710 = ~ ( n33 ) ;
assign n711 =  ( n709 ) & ( n710 )  ;
assign n712 = ~ ( n38 ) ;
assign n713 =  ( n711 ) & ( n712 )  ;
assign n714 = ~ ( n43 ) ;
assign n715 =  ( n713 ) & ( n714 )  ;
assign n716 =  ( n713 ) & ( n43 )  ;
assign n717 =  ( n711 ) & ( n38 )  ;
assign n718 = ~ ( n387 ) ;
assign n719 =  ( n717 ) & ( n718 )  ;
assign n720 =  ( n717 ) & ( n387 )  ;
assign n721 =  ( n709 ) & ( n33 )  ;
assign n722 =  ( n707 ) & ( n24 )  ;
assign n723 =  ( n705 ) & ( n15 )  ;
assign n724 =  ( n703 ) & ( n11 )  ;
assign LB2D_proc_0_addr0 = n720 ? (n388) : (0);
assign LB2D_proc_0_data0 = n720 ? (n386) : (LB2D_proc_0[0]);
assign n725 = ~ ( n390 ) ;
assign n726 =  ( n717 ) & ( n725 )  ;
assign n727 =  ( n717 ) & ( n390 )  ;
assign LB2D_proc_1_addr0 = n727 ? (n388) : (0);
assign LB2D_proc_1_data0 = n727 ? (n386) : (LB2D_proc_1[0]);
assign n728 = ~ ( n392 ) ;
assign n729 =  ( n717 ) & ( n728 )  ;
assign n730 =  ( n717 ) & ( n392 )  ;
assign LB2D_proc_2_addr0 = n730 ? (n388) : (0);
assign LB2D_proc_2_data0 = n730 ? (n386) : (LB2D_proc_2[0]);
assign n731 = ~ ( n394 ) ;
assign n732 =  ( n717 ) & ( n731 )  ;
assign n733 =  ( n717 ) & ( n394 )  ;
assign LB2D_proc_3_addr0 = n733 ? (n388) : (0);
assign LB2D_proc_3_data0 = n733 ? (n386) : (LB2D_proc_3[0]);
assign n734 = ~ ( n396 ) ;
assign n735 =  ( n717 ) & ( n734 )  ;
assign n736 =  ( n717 ) & ( n396 )  ;
assign LB2D_proc_4_addr0 = n736 ? (n388) : (0);
assign LB2D_proc_4_data0 = n736 ? (n386) : (LB2D_proc_4[0]);
assign n737 = ~ ( n398 ) ;
assign n738 =  ( n717 ) & ( n737 )  ;
assign n739 =  ( n717 ) & ( n398 )  ;
assign LB2D_proc_5_addr0 = n739 ? (n388) : (0);
assign LB2D_proc_5_data0 = n739 ? (n386) : (LB2D_proc_5[0]);
assign n740 = ~ ( n400 ) ;
assign n741 =  ( n717 ) & ( n740 )  ;
assign n742 =  ( n717 ) & ( n400 )  ;
assign LB2D_proc_6_addr0 = n742 ? (n388) : (0);
assign LB2D_proc_6_data0 = n742 ? (n386) : (LB2D_proc_6[0]);
assign n743 = ~ ( n80 ) ;
assign n744 =  ( n717 ) & ( n743 )  ;
assign n745 =  ( n717 ) & ( n80 )  ;
assign LB2D_proc_7_addr0 = n745 ? (n388) : (0);
assign LB2D_proc_7_data0 = n745 ? (n386) : (LB2D_proc_7[0]);
/*
function [7:0] gb_fun ;
input [647:0] arg0;
    begin
//TODO: Add the specific function HERE.    end
endfunction
*/

always @(posedge clk) begin
   if(rst) begin
       LB1D_buff <= LB1D_buff;
       LB1D_in <= LB1D_in;
       LB1D_it_1 <= LB1D_it_1;
       LB1D_p_cnt <= LB1D_p_cnt;
       LB1D_uIn <= LB1D_uIn;
       LB2D_proc_w <= LB2D_proc_w;
       LB2D_proc_x <= LB2D_proc_x;
       LB2D_proc_y <= LB2D_proc_y;
       LB2D_shift_0 <= LB2D_shift_0;
       LB2D_shift_1 <= LB2D_shift_1;
       LB2D_shift_2 <= LB2D_shift_2;
       LB2D_shift_3 <= LB2D_shift_3;
       LB2D_shift_4 <= LB2D_shift_4;
       LB2D_shift_5 <= LB2D_shift_5;
       LB2D_shift_6 <= LB2D_shift_6;
       LB2D_shift_7 <= LB2D_shift_7;
       LB2D_shift_x <= LB2D_shift_x;
       LB2D_shift_y <= LB2D_shift_y;
       arg_0_TDATA <= arg_0_TDATA;
       arg_0_TVALID <= arg_0_TVALID;
       arg_1_TREADY <= arg_1_TREADY;
       gb_exit_it_1 <= gb_exit_it_1;
       gb_exit_it_2 <= gb_exit_it_2;
       gb_exit_it_3 <= gb_exit_it_3;
       gb_exit_it_4 <= gb_exit_it_4;
       gb_exit_it_5 <= gb_exit_it_5;
       gb_exit_it_6 <= gb_exit_it_6;
       gb_exit_it_7 <= gb_exit_it_7;
       gb_exit_it_8 <= gb_exit_it_8;
       gb_p_cnt <= gb_p_cnt;
       gb_pp_it_1 <= gb_pp_it_1;
       gb_pp_it_2 <= gb_pp_it_2;
       gb_pp_it_3 <= gb_pp_it_3;
       gb_pp_it_4 <= gb_pp_it_4;
       gb_pp_it_5 <= gb_pp_it_5;
       gb_pp_it_6 <= gb_pp_it_6;
       gb_pp_it_7 <= gb_pp_it_7;
       gb_pp_it_8 <= gb_pp_it_8;
       gb_pp_it_9 <= gb_pp_it_9;
       in_stream_buff_0 <= in_stream_buff_0;
       in_stream_buff_1 <= in_stream_buff_1;
       in_stream_empty <= in_stream_empty;
       in_stream_full <= in_stream_full;
       slice_stream_buff_0 <= slice_stream_buff_0;
       slice_stream_buff_1 <= slice_stream_buff_1;
       slice_stream_empty <= slice_stream_empty;
       slice_stream_full <= slice_stream_full;
       stencil_stream_buff_0 <= stencil_stream_buff_0;
       stencil_stream_buff_1 <= stencil_stream_buff_1;
       stencil_stream_empty <= stencil_stream_empty;
       stencil_stream_full <= stencil_stream_full;
   end
   else if(step) begin
       LB1D_buff <= n51;
       LB1D_in <= n59;
       LB1D_it_1 <= n62;
       LB1D_p_cnt <= n71;
       LB1D_uIn <= n78;
       LB2D_proc_w <= n90;
       LB2D_proc_x <= n99;
       LB2D_proc_y <= n110;
       LB2D_shift_0 <= n117;
       LB2D_shift_1 <= n124;
       LB2D_shift_2 <= n131;
       LB2D_shift_3 <= n138;
       LB2D_shift_4 <= n145;
       LB2D_shift_5 <= n152;
       LB2D_shift_6 <= n159;
       LB2D_shift_7 <= n168;
       LB2D_shift_x <= n181;
       LB2D_shift_y <= n193;
       arg_0_TDATA <= n203;
       arg_0_TVALID <= n214;
       arg_1_TREADY <= n222;
       gb_exit_it_1 <= n231;
       gb_exit_it_2 <= n238;
       gb_exit_it_3 <= n245;
       gb_exit_it_4 <= n252;
       gb_exit_it_5 <= n259;
       gb_exit_it_6 <= n266;
       gb_exit_it_7 <= n273;
       gb_exit_it_8 <= n280;
       gb_p_cnt <= n290;
       gb_pp_it_1 <= n297;
       gb_pp_it_2 <= n304;
       gb_pp_it_3 <= n311;
       gb_pp_it_4 <= n318;
       gb_pp_it_5 <= n325;
       gb_pp_it_6 <= n332;
       gb_pp_it_7 <= n339;
       gb_pp_it_8 <= n346;
       gb_pp_it_9 <= n353;
       in_stream_buff_0 <= n360;
       in_stream_buff_1 <= n367;
       in_stream_empty <= n376;
       in_stream_full <= n385;
       slice_stream_buff_0 <= n474;
       slice_stream_buff_1 <= n482;
       slice_stream_empty <= n491;
       slice_stream_full <= n501;
       stencil_stream_buff_0 <= n673;
       stencil_stream_buff_1 <= n681;
       stencil_stream_empty <= n691;
       stencil_stream_full <= n702;
       LB2D_proc_0 [ LB2D_proc_0_addr0 ] <= LB2D_proc_0_data0;
       LB2D_proc_1 [ LB2D_proc_1_addr0 ] <= LB2D_proc_1_data0;
       LB2D_proc_2 [ LB2D_proc_2_addr0 ] <= LB2D_proc_2_data0;
       LB2D_proc_3 [ LB2D_proc_3_addr0 ] <= LB2D_proc_3_data0;
       LB2D_proc_4 [ LB2D_proc_4_addr0 ] <= LB2D_proc_4_data0;
       LB2D_proc_5 [ LB2D_proc_5_addr0 ] <= LB2D_proc_5_data0;
       LB2D_proc_6 [ LB2D_proc_6_addr0 ] <= LB2D_proc_6_data0;
       LB2D_proc_7 [ LB2D_proc_7_addr0 ] <= LB2D_proc_7_data0;
   end
end
endmodule
