module SPEC_B(
arg_0_TREADY,
arg_1_TDATA,
arg_1_TVALID,
LB1D_buff,
LB1D_in,
LB1D_it_1,
LB1D_p_cnt,
LB1D_uIn,
LB2D_proc_w,
LB2D_proc_x,
LB2D_proc_y,
LB2D_shift_0,
LB2D_shift_1,
LB2D_shift_2,
LB2D_shift_3,
LB2D_shift_4,
LB2D_shift_5,
LB2D_shift_6,
LB2D_shift_7,
LB2D_shift_x,
LB2D_shift_y,
arg_0_TDATA,
arg_0_TVALID,
arg_1_TREADY,
gb_exit_it_1,
gb_exit_it_2,
gb_exit_it_3,
gb_exit_it_4,
gb_exit_it_5,
gb_exit_it_6,
gb_exit_it_7,
gb_exit_it_8,
gb_p_cnt,
gb_pp_it_1,
gb_pp_it_2,
gb_pp_it_3,
gb_pp_it_4,
gb_pp_it_5,
gb_pp_it_6,
gb_pp_it_7,
gb_pp_it_8,
gb_pp_it_9,
in_stream_buff_0,
in_stream_buff_1,
in_stream_empty,
in_stream_full,
slice_stream_buff_0,
slice_stream_buff_1,
slice_stream_empty,
slice_stream_full,
stencil_stream_buff_0,
stencil_stream_buff_1,
stencil_stream_empty,
stencil_stream_full,
clk,rst,
step
);
input            arg_0_TREADY;
input      [7:0] arg_1_TDATA;
input            arg_1_TVALID;
input clk;
input rst;
input step;
output      [7:0] LB1D_buff;
output      [7:0] LB1D_in;
output            LB1D_it_1;
output     [18:0] LB1D_p_cnt;
output      [7:0] LB1D_uIn;
output     [63:0] LB2D_proc_w;
output      [8:0] LB2D_proc_x;
output      [9:0] LB2D_proc_y;
output     [71:0] LB2D_shift_0;
output     [71:0] LB2D_shift_1;
output     [71:0] LB2D_shift_2;
output     [71:0] LB2D_shift_3;
output     [71:0] LB2D_shift_4;
output     [71:0] LB2D_shift_5;
output     [71:0] LB2D_shift_6;
output     [71:0] LB2D_shift_7;
output      [8:0] LB2D_shift_x;
output      [9:0] LB2D_shift_y;
output      [7:0] arg_0_TDATA;
output            arg_0_TVALID;
output            arg_1_TREADY;
output            gb_exit_it_1;
output            gb_exit_it_2;
output            gb_exit_it_3;
output            gb_exit_it_4;
output            gb_exit_it_5;
output            gb_exit_it_6;
output            gb_exit_it_7;
output            gb_exit_it_8;
output     [18:0] gb_p_cnt;
output            gb_pp_it_1;
output            gb_pp_it_2;
output            gb_pp_it_3;
output            gb_pp_it_4;
output            gb_pp_it_5;
output            gb_pp_it_6;
output            gb_pp_it_7;
output            gb_pp_it_8;
output            gb_pp_it_9;
output      [7:0] in_stream_buff_0;
output      [7:0] in_stream_buff_1;
output            in_stream_empty;
output            in_stream_full;
output     [71:0] slice_stream_buff_0;
output     [71:0] slice_stream_buff_1;
output            slice_stream_empty;
output            slice_stream_full;
output    [647:0] stencil_stream_buff_0;
output    [647:0] stencil_stream_buff_1;
output            stencil_stream_empty;
output            stencil_stream_full;
reg      [7:0] LB1D_buff;
reg      [7:0] LB1D_in;
reg            LB1D_it_1;
reg     [18:0] LB1D_p_cnt;
reg      [7:0] LB1D_uIn;
reg     [63:0] LB2D_proc_w;
reg      [8:0] LB2D_proc_x;
reg      [9:0] LB2D_proc_y;
reg     [71:0] LB2D_shift_0;
reg     [71:0] LB2D_shift_1;
reg     [71:0] LB2D_shift_2;
reg     [71:0] LB2D_shift_3;
reg     [71:0] LB2D_shift_4;
reg     [71:0] LB2D_shift_5;
reg     [71:0] LB2D_shift_6;
reg     [71:0] LB2D_shift_7;
reg      [8:0] LB2D_shift_x;
reg      [9:0] LB2D_shift_y;
reg      [7:0] arg_0_TDATA;
reg            arg_0_TVALID;
reg            arg_1_TREADY;
reg            gb_exit_it_1;
reg            gb_exit_it_2;
reg            gb_exit_it_3;
reg            gb_exit_it_4;
reg            gb_exit_it_5;
reg            gb_exit_it_6;
reg            gb_exit_it_7;
reg            gb_exit_it_8;
reg     [18:0] gb_p_cnt;
reg            gb_pp_it_1;
reg            gb_pp_it_2;
reg            gb_pp_it_3;
reg            gb_pp_it_4;
reg            gb_pp_it_5;
reg            gb_pp_it_6;
reg            gb_pp_it_7;
reg            gb_pp_it_8;
reg            gb_pp_it_9;
reg      [7:0] in_stream_buff_0;
reg      [7:0] in_stream_buff_1;
reg            in_stream_empty;
reg            in_stream_full;
reg     [71:0] slice_stream_buff_0;
reg     [71:0] slice_stream_buff_1;
reg            slice_stream_empty;
reg            slice_stream_full;
reg    [647:0] stencil_stream_buff_0;
reg    [647:0] stencil_stream_buff_1;
reg            stencil_stream_empty;
reg            stencil_stream_full;
wire            arg_0_TREADY;
wire      [7:0] arg_1_TDATA;
wire            arg_1_TVALID;
wire            n0;
wire            n1;
wire            n2;
wire            n3;
wire            n4;
wire            n5;
wire            n6;
wire            n7;
wire            n8;
wire            n9;
wire            n10;
wire            n11;
wire            n12;
wire            n13;
wire            n14;
wire            n15;
wire            n16;
wire            n17;
wire            n18;
wire            n19;
wire            n20;
wire            n21;
wire            n22;
wire            n23;
wire            n24;
wire            n25;
wire            n26;
wire            n27;
wire            n28;
wire            n29;
wire            n30;
wire            n31;
wire            n32;
wire            n33;
wire            n34;
wire      [7:0] n35;
wire      [7:0] n36;
wire      [7:0] n37;
wire      [7:0] n38;
wire      [7:0] n39;
wire      [7:0] n40;
wire      [7:0] n41;
wire      [7:0] n42;
wire      [7:0] n43;
wire      [7:0] n44;
wire      [7:0] n45;
wire      [7:0] n46;
wire            n47;
wire            n48;
wire            n49;
wire            n50;
wire     [18:0] n51;
wire     [18:0] n52;
wire     [18:0] n53;
wire     [18:0] n54;
wire     [18:0] n55;
wire     [18:0] n56;
wire     [18:0] n57;
wire     [18:0] n58;
wire      [7:0] n59;
wire      [7:0] n60;
wire      [7:0] n61;
wire      [7:0] n62;
wire      [7:0] n63;
wire            n64;
wire            n65;
wire     [63:0] n66;
wire     [63:0] n67;
wire     [63:0] n68;
wire     [63:0] n69;
wire     [63:0] n70;
wire     [63:0] n71;
wire     [63:0] n72;
wire     [63:0] n73;
wire      [8:0] n74;
wire      [8:0] n75;
wire      [8:0] n76;
wire      [8:0] n77;
wire      [8:0] n78;
wire      [8:0] n79;
wire      [8:0] n80;
wire            n81;
wire      [9:0] n82;
wire      [9:0] n83;
wire      [9:0] n84;
wire      [9:0] n85;
wire      [9:0] n86;
wire      [9:0] n87;
wire      [9:0] n88;
wire      [9:0] n89;
wire     [71:0] n90;
wire     [71:0] n91;
wire     [71:0] n92;
wire     [71:0] n93;
wire     [71:0] n94;
wire     [71:0] n95;
wire     [71:0] n96;
wire     [71:0] n97;
wire     [71:0] n98;
wire     [71:0] n99;
wire     [71:0] n100;
wire     [71:0] n101;
wire     [71:0] n102;
wire     [71:0] n103;
wire     [71:0] n104;
wire     [71:0] n105;
wire     [71:0] n106;
wire     [71:0] n107;
wire     [71:0] n108;
wire     [71:0] n109;
wire     [71:0] n110;
wire     [71:0] n111;
wire     [71:0] n112;
wire     [71:0] n113;
wire     [71:0] n114;
wire     [71:0] n115;
wire     [71:0] n116;
wire     [71:0] n117;
wire     [71:0] n118;
wire     [71:0] n119;
wire     [71:0] n120;
wire     [71:0] n121;
wire     [71:0] n122;
wire     [71:0] n123;
wire     [71:0] n124;
wire            n125;
wire     [71:0] n126;
wire     [71:0] n127;
wire     [71:0] n128;
wire     [71:0] n129;
wire     [71:0] n130;
wire     [71:0] n131;
wire      [8:0] n132;
wire      [8:0] n133;
wire      [8:0] n134;
wire      [8:0] n135;
wire      [8:0] n136;
wire      [8:0] n137;
wire            n138;
wire            n139;
wire      [9:0] n140;
wire      [9:0] n141;
wire      [9:0] n142;
wire      [9:0] n143;
wire      [9:0] n144;
wire      [9:0] n145;
wire      [9:0] n146;
wire      [9:0] n147;
wire            n148;
wire    [647:0] n149;
wire      [7:0] n150;
wire      [7:0] n151;
wire      [7:0] n152;
wire      [7:0] n153;
wire      [7:0] n154;
wire      [7:0] n155;
wire            n156;
wire            n157;
wire            n158;
wire            n159;
wire            n160;
wire            n161;
wire            n162;
wire     [18:0] n163;
wire            n164;
wire            n165;
wire            n166;
wire            n167;
wire            n168;
wire            n169;
wire            n170;
wire            n171;
wire     [18:0] n172;
wire            n173;
wire            n174;
wire            n175;
wire            n176;
wire            n177;
wire            n178;
wire            n179;
wire            n180;
wire            n181;
wire            n182;
wire            n183;
wire            n184;
wire            n185;
wire            n186;
wire            n187;
wire            n188;
wire            n189;
wire            n190;
wire            n191;
wire            n192;
wire            n193;
wire            n194;
wire            n195;
wire            n196;
wire            n197;
wire            n198;
wire            n199;
wire            n200;
wire            n201;
wire            n202;
wire            n203;
wire            n204;
wire            n205;
wire            n206;
wire            n207;
wire            n208;
wire            n209;
wire            n210;
wire            n211;
wire            n212;
wire            n213;
wire            n214;
wire            n215;
wire     [18:0] n216;
wire     [18:0] n217;
wire     [18:0] n218;
wire     [18:0] n219;
wire     [18:0] n220;
wire     [18:0] n221;
wire            n222;
wire            n223;
wire            n224;
wire            n225;
wire            n226;
wire            n227;
wire            n228;
wire            n229;
wire            n230;
wire            n231;
wire            n232;
wire            n233;
wire            n234;
wire            n235;
wire            n236;
wire            n237;
wire            n238;
wire            n239;
wire            n240;
wire            n241;
wire            n242;
wire            n243;
wire            n244;
wire            n245;
wire            n246;
wire            n247;
wire            n248;
wire            n249;
wire            n250;
wire            n251;
wire            n252;
wire            n253;
wire            n254;
wire            n255;
wire            n256;
wire            n257;
wire            n258;
wire            n259;
wire            n260;
wire            n261;
wire            n262;
wire            n263;
wire            n264;
wire            n265;
wire            n266;
wire      [7:0] n267;
wire      [7:0] n268;
wire      [7:0] n269;
wire      [7:0] n270;
wire      [7:0] n271;
wire      [7:0] n272;
wire      [7:0] n273;
wire      [7:0] n274;
wire      [7:0] n275;
wire      [7:0] n276;
wire            n277;
wire            n278;
wire            n279;
wire            n280;
wire            n281;
wire            n282;
wire            n283;
wire            n284;
wire            n285;
wire            n286;
wire            n287;
wire            n288;
wire            n289;
wire            n290;
wire      [7:0] n291;
wire            n292;
wire      [8:0] n293;
wire      [7:0] n294;
wire            n295;
wire      [7:0] n296;
wire            n297;
wire      [7:0] n298;
wire            n299;
wire      [7:0] n300;
wire            n301;
wire      [7:0] n302;
wire            n303;
wire      [7:0] n304;
wire            n305;
wire      [7:0] n306;
wire      [7:0] n307;
wire      [7:0] n308;
wire      [7:0] n309;
wire      [7:0] n310;
wire      [7:0] n311;
wire      [7:0] n312;
wire      [7:0] n313;
wire      [7:0] n314;
wire      [7:0] n315;
wire      [7:0] n316;
wire      [7:0] n317;
wire      [7:0] n318;
wire      [7:0] n319;
wire      [7:0] n320;
wire      [7:0] n321;
wire      [7:0] n322;
wire      [7:0] n323;
wire      [7:0] n324;
wire      [7:0] n325;
wire      [7:0] n326;
wire      [7:0] n327;
wire      [7:0] n328;
wire      [7:0] n329;
wire      [7:0] n330;
wire      [7:0] n331;
wire      [7:0] n332;
wire      [7:0] n333;
wire      [7:0] n334;
wire      [7:0] n335;
wire      [7:0] n336;
wire      [7:0] n337;
wire      [7:0] n338;
wire      [7:0] n339;
wire      [7:0] n340;
wire      [7:0] n341;
wire      [7:0] n342;
wire      [7:0] n343;
wire      [7:0] n344;
wire      [7:0] n345;
wire      [7:0] n346;
wire      [7:0] n347;
wire      [7:0] n348;
wire      [7:0] n349;
wire      [7:0] n350;
wire      [7:0] n351;
wire      [7:0] n352;
wire      [7:0] n353;
wire      [7:0] n354;
wire      [7:0] n355;
wire      [7:0] n356;
wire      [7:0] n357;
wire      [7:0] n358;
wire      [7:0] n359;
wire      [7:0] n360;
wire      [7:0] n361;
wire      [7:0] n362;
wire      [7:0] n363;
wire     [15:0] n364;
wire     [23:0] n365;
wire     [31:0] n366;
wire     [39:0] n367;
wire     [47:0] n368;
wire     [55:0] n369;
wire     [63:0] n370;
wire     [71:0] n371;
wire     [71:0] n372;
wire     [71:0] n373;
wire     [71:0] n374;
wire     [71:0] n375;
wire     [71:0] n376;
wire     [71:0] n377;
wire     [71:0] n378;
wire     [71:0] n379;
wire     [71:0] n380;
wire     [71:0] n381;
wire     [71:0] n382;
wire     [71:0] n383;
wire            n384;
wire            n385;
wire            n386;
wire            n387;
wire            n388;
wire            n389;
wire            n390;
wire            n391;
wire            n392;
wire            n393;
wire            n394;
wire            n395;
wire            n396;
wire            n397;
wire            n398;
wire            n399;
wire            n400;
wire            n401;
wire      [7:0] n402;
wire      [7:0] n403;
wire      [7:0] n404;
wire      [7:0] n405;
wire      [7:0] n406;
wire      [7:0] n407;
wire      [7:0] n408;
wire      [7:0] n409;
wire      [7:0] n410;
wire     [15:0] n411;
wire     [23:0] n412;
wire     [31:0] n413;
wire     [39:0] n414;
wire     [47:0] n415;
wire     [55:0] n416;
wire     [63:0] n417;
wire     [71:0] n418;
wire      [7:0] n419;
wire      [7:0] n420;
wire      [7:0] n421;
wire      [7:0] n422;
wire      [7:0] n423;
wire      [7:0] n424;
wire      [7:0] n425;
wire      [7:0] n426;
wire      [7:0] n427;
wire     [15:0] n428;
wire     [23:0] n429;
wire     [31:0] n430;
wire     [39:0] n431;
wire     [47:0] n432;
wire     [55:0] n433;
wire     [63:0] n434;
wire     [71:0] n435;
wire      [7:0] n436;
wire      [7:0] n437;
wire      [7:0] n438;
wire      [7:0] n439;
wire      [7:0] n440;
wire      [7:0] n441;
wire      [7:0] n442;
wire      [7:0] n443;
wire      [7:0] n444;
wire     [15:0] n445;
wire     [23:0] n446;
wire     [31:0] n447;
wire     [39:0] n448;
wire     [47:0] n449;
wire     [55:0] n450;
wire     [63:0] n451;
wire     [71:0] n452;
wire      [7:0] n453;
wire      [7:0] n454;
wire      [7:0] n455;
wire      [7:0] n456;
wire      [7:0] n457;
wire      [7:0] n458;
wire      [7:0] n459;
wire      [7:0] n460;
wire      [7:0] n461;
wire     [15:0] n462;
wire     [23:0] n463;
wire     [31:0] n464;
wire     [39:0] n465;
wire     [47:0] n466;
wire     [55:0] n467;
wire     [63:0] n468;
wire     [71:0] n469;
wire      [7:0] n470;
wire      [7:0] n471;
wire      [7:0] n472;
wire      [7:0] n473;
wire      [7:0] n474;
wire      [7:0] n475;
wire      [7:0] n476;
wire      [7:0] n477;
wire      [7:0] n478;
wire     [15:0] n479;
wire     [23:0] n480;
wire     [31:0] n481;
wire     [39:0] n482;
wire     [47:0] n483;
wire     [55:0] n484;
wire     [63:0] n485;
wire     [71:0] n486;
wire      [7:0] n487;
wire      [7:0] n488;
wire      [7:0] n489;
wire      [7:0] n490;
wire      [7:0] n491;
wire      [7:0] n492;
wire      [7:0] n493;
wire      [7:0] n494;
wire      [7:0] n495;
wire     [15:0] n496;
wire     [23:0] n497;
wire     [31:0] n498;
wire     [39:0] n499;
wire     [47:0] n500;
wire     [55:0] n501;
wire     [63:0] n502;
wire     [71:0] n503;
wire      [7:0] n504;
wire      [7:0] n505;
wire      [7:0] n506;
wire      [7:0] n507;
wire      [7:0] n508;
wire      [7:0] n509;
wire      [7:0] n510;
wire      [7:0] n511;
wire      [7:0] n512;
wire     [15:0] n513;
wire     [23:0] n514;
wire     [31:0] n515;
wire     [39:0] n516;
wire     [47:0] n517;
wire     [55:0] n518;
wire     [63:0] n519;
wire     [71:0] n520;
wire      [7:0] n521;
wire      [7:0] n522;
wire      [7:0] n523;
wire      [7:0] n524;
wire      [7:0] n525;
wire      [7:0] n526;
wire      [7:0] n527;
wire      [7:0] n528;
wire      [7:0] n529;
wire     [15:0] n530;
wire     [23:0] n531;
wire     [31:0] n532;
wire     [39:0] n533;
wire     [47:0] n534;
wire     [55:0] n535;
wire     [63:0] n536;
wire     [71:0] n537;
wire      [7:0] n538;
wire      [7:0] n539;
wire      [7:0] n540;
wire      [7:0] n541;
wire      [7:0] n542;
wire      [7:0] n543;
wire      [7:0] n544;
wire      [7:0] n545;
wire      [7:0] n546;
wire     [15:0] n547;
wire     [23:0] n548;
wire     [31:0] n549;
wire     [39:0] n550;
wire     [47:0] n551;
wire     [55:0] n552;
wire     [63:0] n553;
wire     [71:0] n554;
wire    [143:0] n555;
wire    [215:0] n556;
wire    [287:0] n557;
wire    [359:0] n558;
wire    [431:0] n559;
wire    [503:0] n560;
wire    [575:0] n561;
wire    [647:0] n562;
wire    [647:0] n563;
wire    [647:0] n564;
wire    [647:0] n565;
wire    [647:0] n566;
wire    [647:0] n567;
wire    [647:0] n568;
wire    [647:0] n569;
wire    [647:0] n570;
wire    [647:0] n571;
wire    [647:0] n572;
wire    [647:0] n573;
wire            n574;
wire            n575;
wire            n576;
wire            n577;
wire            n578;
wire            n579;
wire            n580;
wire            n581;
wire            n582;
wire            n583;
wire            n584;
wire            n585;
wire            n586;
wire            n587;
wire            n588;
wire            n589;
wire            n590;
wire      [8:0] LB2D_proc_0_addr0;
wire      [7:0] LB2D_proc_0_data0;
wire            n591;
wire            n592;
wire            n593;
wire            n594;
wire            n595;
wire            n596;
wire            n597;
wire            n598;
wire            n599;
wire            n600;
wire            n601;
wire            n602;
wire            n603;
wire            n604;
wire            n605;
wire            n606;
wire      [8:0] LB2D_proc_1_addr0;
wire      [7:0] LB2D_proc_1_data0;
wire            n607;
wire            n608;
wire            n609;
wire      [8:0] LB2D_proc_2_addr0;
wire      [7:0] LB2D_proc_2_data0;
wire            n610;
wire            n611;
wire            n612;
wire      [8:0] LB2D_proc_3_addr0;
wire      [7:0] LB2D_proc_3_data0;
wire            n613;
wire            n614;
wire            n615;
wire      [8:0] LB2D_proc_4_addr0;
wire      [7:0] LB2D_proc_4_data0;
wire            n616;
wire            n617;
wire            n618;
wire      [8:0] LB2D_proc_5_addr0;
wire      [7:0] LB2D_proc_5_data0;
wire            n619;
wire            n620;
wire            n621;
wire      [8:0] LB2D_proc_6_addr0;
wire      [7:0] LB2D_proc_6_data0;
wire            n622;
wire            n623;
wire            n624;
wire      [8:0] LB2D_proc_7_addr0;
wire      [7:0] LB2D_proc_7_data0;
wire            n625;
wire            n626;
wire            n627;
reg      [7:0] LB2D_proc_0[487:0];
reg      [7:0] LB2D_proc_1[487:0];
reg      [7:0] LB2D_proc_2[487:0];
reg      [7:0] LB2D_proc_3[487:0];
reg      [7:0] LB2D_proc_4[487:0];
reg      [7:0] LB2D_proc_5[487:0];
reg      [7:0] LB2D_proc_6[487:0];
reg      [7:0] LB2D_proc_7[487:0];
wire clk;
wire rst;
wire step;
assign n0 =  ( arg_0_TREADY ) == ( 1'd1 )  ;
assign n1 =  ( arg_0_TVALID ) == ( 1'd1 )  ;
assign n2 =  ( n0 ) & ( n1 )  ;
assign n3 =  ( arg_1_TVALID ) == ( 1'd0 )  ;
assign n4 =  ( n2 ) & ( n3 )  ;
assign n5 =  ( arg_0_TVALID ) == ( 1'd0 )  ;
assign n6 =  ( gb_exit_it_1 ) == ( 1'd0 )  ;
assign n7 =  ( stencil_stream_empty ) == ( 1'd0 )  ;
assign n8 =  ( n6 ) & ( n7 )  ;
assign n9 =  ( gb_exit_it_1 ) == ( 1'd1 )  ;
assign n10 =  ( gb_exit_it_8 ) == ( 1'd0 )  ;
assign n11 =  ( n9 ) & ( n10 )  ;
assign n12 =  ( n8 ) | ( n11 )  ;
assign n13 =  ( n5 ) & ( n12 )  ;
assign n14 =  ( slice_stream_empty ) == ( 1'd0 )  ;
assign n15 =  ( LB2D_shift_x ) != ( 9'd488 )  ;
assign n16 =  ( n14 ) & ( n15 )  ;
assign n17 =  ( stencil_stream_full ) == ( 1'd0 )  ;
assign n18 =  ( LB2D_shift_x ) < ( 9'd8 )  ;
assign n19 =  ( LB2D_shift_x ) > ( 9'd0 )  ;
assign n20 =  ( n18 ) & ( n19 )  ;
assign n21 =  ( n17 ) | ( n20 )  ;
assign n22 =  ( n16 ) & ( n21 )  ;
assign n23 =  ( in_stream_empty ) == ( 1'd0 )  ;
assign n24 =  ( slice_stream_full ) == ( 1'd0 )  ;
assign n25 =  ( LB2D_proc_y ) < ( 10'd8 )  ;
assign n26 =  ( n24 ) | ( n25 )  ;
assign n27 =  ( n23 ) & ( n26 )  ;
assign n28 =  ( arg_1_TREADY ) == ( 1'd0 )  ;
assign n29 =  ( in_stream_full ) == ( 1'd0 )  ;
assign n30 =  ( n28 ) & ( n29 )  ;
assign n31 =  ( LB1D_it_1 ) == ( 1'd0 )  ;
assign n32 =  ( n30 ) & ( n31 )  ;
assign n33 =  ( LB1D_it_1 ) == ( 1'd1 )  ;
assign n34 =  ( n30 ) & ( n33 )  ;
assign n35 =  ( n34 ) ? ( LB1D_uIn ) : ( LB1D_buff ) ;
assign n36 =  ( n32 ) ? ( LB1D_uIn ) : ( n35 ) ;
assign n37 =  ( n27 ) ? ( LB1D_buff ) : ( n36 ) ;
assign n38 =  ( n22 ) ? ( LB1D_buff ) : ( n37 ) ;
assign n39 =  ( n13 ) ? ( LB1D_buff ) : ( n38 ) ;
assign n40 =  ( n4 ) ? ( LB1D_buff ) : ( n39 ) ;
assign n41 =  ( n34 ) ? ( LB1D_in ) : ( LB1D_in ) ;
assign n42 =  ( n32 ) ? ( LB1D_in ) : ( n41 ) ;
assign n43 =  ( n27 ) ? ( LB1D_in ) : ( n42 ) ;
assign n44 =  ( n22 ) ? ( LB1D_in ) : ( n43 ) ;
assign n45 =  ( n13 ) ? ( LB1D_in ) : ( n44 ) ;
assign n46 =  ( n4 ) ? ( LB1D_in ) : ( n45 ) ;
assign n47 =  ( LB1D_p_cnt ) == ( 19'd316224 )  ;
assign n48 =  ( n47 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n49 =  ( n34 ) ? ( n48 ) : ( LB1D_it_1 ) ;
assign n50 =  ( n32 ) ? ( 1'd1 ) : ( n49 ) ;
assign n51 =  ( LB1D_p_cnt ) + ( 19'd1 )  ;
assign n52 =  ( n47 ) ? ( 19'd0 ) : ( n51 ) ;
assign n53 =  ( n34 ) ? ( n52 ) : ( LB1D_p_cnt ) ;
assign n54 =  ( n32 ) ? ( n51 ) : ( n53 ) ;
assign n55 =  ( n27 ) ? ( LB1D_p_cnt ) : ( n54 ) ;
assign n56 =  ( n22 ) ? ( LB1D_p_cnt ) : ( n55 ) ;
assign n57 =  ( n13 ) ? ( LB1D_p_cnt ) : ( n56 ) ;
assign n58 =  ( n4 ) ? ( LB1D_p_cnt ) : ( n57 ) ;
assign n59 =  ( n34 ) ? ( LB1D_in ) : ( LB1D_uIn ) ;
assign n60 =  ( n32 ) ? ( LB1D_in ) : ( n59 ) ;
assign n61 =  ( n27 ) ? ( LB1D_uIn ) : ( n60 ) ;
assign n62 =  ( n22 ) ? ( LB1D_uIn ) : ( n61 ) ;
assign n63 =  ( n13 ) ? ( LB1D_uIn ) : ( n62 ) ;
assign n64 =  ( LB2D_proc_x ) == ( 9'd488 )  ;
assign n65 =  ( LB2D_proc_w ) == ( 64'd7 )  ;
assign n66 =  ( LB2D_proc_w ) + ( 64'd1 )  ;
assign n67 =  ( n65 ) ? ( 64'd0 ) : ( n66 ) ;
assign n68 =  ( n64 ) ? ( n67 ) : ( LB2D_proc_w ) ;
assign n69 =  ( n34 ) ? ( LB2D_proc_w ) : ( LB2D_proc_w ) ;
assign n70 =  ( n27 ) ? ( n68 ) : ( n69 ) ;
assign n71 =  ( n22 ) ? ( LB2D_proc_w ) : ( n70 ) ;
assign n72 =  ( n13 ) ? ( LB2D_proc_w ) : ( n71 ) ;
assign n73 =  ( n4 ) ? ( LB2D_proc_w ) : ( n72 ) ;
assign n74 =  ( LB2D_proc_x ) + ( 9'd1 )  ;
assign n75 =  ( n64 ) ? ( 9'd1 ) : ( n74 ) ;
assign n76 =  ( n34 ) ? ( LB2D_proc_x ) : ( LB2D_proc_x ) ;
assign n77 =  ( n27 ) ? ( n75 ) : ( n76 ) ;
assign n78 =  ( n22 ) ? ( LB2D_proc_x ) : ( n77 ) ;
assign n79 =  ( n13 ) ? ( LB2D_proc_x ) : ( n78 ) ;
assign n80 =  ( n4 ) ? ( LB2D_proc_x ) : ( n79 ) ;
assign n81 =  ( LB2D_proc_y ) == ( 10'd648 )  ;
assign n82 =  ( LB2D_proc_y ) + ( 10'd1 )  ;
assign n83 =  ( n81 ) ? ( 10'd0 ) : ( n82 ) ;
assign n84 =  ( n64 ) ? ( n83 ) : ( LB2D_proc_y ) ;
assign n85 =  ( n34 ) ? ( LB2D_proc_y ) : ( LB2D_proc_y ) ;
assign n86 =  ( n27 ) ? ( n84 ) : ( n85 ) ;
assign n87 =  ( n22 ) ? ( LB2D_proc_y ) : ( n86 ) ;
assign n88 =  ( n13 ) ? ( LB2D_proc_y ) : ( n87 ) ;
assign n89 =  ( n4 ) ? ( LB2D_proc_y ) : ( n88 ) ;
assign n90 =  ( n34 ) ? ( LB2D_shift_0 ) : ( LB2D_shift_0 ) ;
assign n91 =  ( n27 ) ? ( LB2D_shift_0 ) : ( n90 ) ;
assign n92 =  ( n22 ) ? ( LB2D_shift_1 ) : ( n91 ) ;
assign n93 =  ( n13 ) ? ( LB2D_shift_0 ) : ( n92 ) ;
assign n94 =  ( n4 ) ? ( LB2D_shift_0 ) : ( n93 ) ;
assign n95 =  ( n34 ) ? ( LB2D_shift_1 ) : ( LB2D_shift_1 ) ;
assign n96 =  ( n27 ) ? ( LB2D_shift_1 ) : ( n95 ) ;
assign n97 =  ( n22 ) ? ( LB2D_shift_2 ) : ( n96 ) ;
assign n98 =  ( n13 ) ? ( LB2D_shift_1 ) : ( n97 ) ;
assign n99 =  ( n4 ) ? ( LB2D_shift_1 ) : ( n98 ) ;
assign n100 =  ( n34 ) ? ( LB2D_shift_2 ) : ( LB2D_shift_2 ) ;
assign n101 =  ( n27 ) ? ( LB2D_shift_2 ) : ( n100 ) ;
assign n102 =  ( n22 ) ? ( LB2D_shift_3 ) : ( n101 ) ;
assign n103 =  ( n13 ) ? ( LB2D_shift_2 ) : ( n102 ) ;
assign n104 =  ( n4 ) ? ( LB2D_shift_2 ) : ( n103 ) ;
assign n105 =  ( n34 ) ? ( LB2D_shift_3 ) : ( LB2D_shift_3 ) ;
assign n106 =  ( n27 ) ? ( LB2D_shift_3 ) : ( n105 ) ;
assign n107 =  ( n22 ) ? ( LB2D_shift_4 ) : ( n106 ) ;
assign n108 =  ( n13 ) ? ( LB2D_shift_3 ) : ( n107 ) ;
assign n109 =  ( n4 ) ? ( LB2D_shift_3 ) : ( n108 ) ;
assign n110 =  ( n34 ) ? ( LB2D_shift_4 ) : ( LB2D_shift_4 ) ;
assign n111 =  ( n27 ) ? ( LB2D_shift_4 ) : ( n110 ) ;
assign n112 =  ( n22 ) ? ( LB2D_shift_5 ) : ( n111 ) ;
assign n113 =  ( n13 ) ? ( LB2D_shift_4 ) : ( n112 ) ;
assign n114 =  ( n4 ) ? ( LB2D_shift_4 ) : ( n113 ) ;
assign n115 =  ( n34 ) ? ( LB2D_shift_5 ) : ( LB2D_shift_5 ) ;
assign n116 =  ( n27 ) ? ( LB2D_shift_5 ) : ( n115 ) ;
assign n117 =  ( n22 ) ? ( LB2D_shift_6 ) : ( n116 ) ;
assign n118 =  ( n13 ) ? ( LB2D_shift_5 ) : ( n117 ) ;
assign n119 =  ( n4 ) ? ( LB2D_shift_5 ) : ( n118 ) ;
assign n120 =  ( n34 ) ? ( LB2D_shift_6 ) : ( LB2D_shift_6 ) ;
assign n121 =  ( n27 ) ? ( LB2D_shift_6 ) : ( n120 ) ;
assign n122 =  ( n22 ) ? ( LB2D_shift_7 ) : ( n121 ) ;
assign n123 =  ( n13 ) ? ( LB2D_shift_6 ) : ( n122 ) ;
assign n124 =  ( n4 ) ? ( LB2D_shift_6 ) : ( n123 ) ;
assign n125 =  ( slice_stream_full ) == ( 1'd1 )  ;
assign n126 =  ( n125 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n127 =  ( n34 ) ? ( LB2D_shift_7 ) : ( LB2D_shift_7 ) ;
assign n128 =  ( n27 ) ? ( LB2D_shift_7 ) : ( n127 ) ;
assign n129 =  ( n22 ) ? ( n126 ) : ( n128 ) ;
assign n130 =  ( n13 ) ? ( LB2D_shift_7 ) : ( n129 ) ;
assign n131 =  ( n4 ) ? ( LB2D_shift_7 ) : ( n130 ) ;
assign n132 =  ( LB2D_shift_x ) + ( 9'd1 )  ;
assign n133 =  ( n34 ) ? ( LB2D_shift_x ) : ( LB2D_shift_x ) ;
assign n134 =  ( n27 ) ? ( LB2D_shift_x ) : ( n133 ) ;
assign n135 =  ( n22 ) ? ( n132 ) : ( n134 ) ;
assign n136 =  ( n13 ) ? ( LB2D_shift_x ) : ( n135 ) ;
assign n137 =  ( n4 ) ? ( LB2D_shift_x ) : ( n136 ) ;
assign n138 =  ( LB2D_shift_y ) < ( 10'd640 )  ;
assign n139 =  ( LB2D_shift_x ) < ( 9'd488 )  ;
assign n140 =  ( LB2D_shift_y ) + ( 10'd1 )  ;
assign n141 =  ( n139 ) ? ( LB2D_shift_y ) : ( n140 ) ;
assign n142 =  ( n138 ) ? ( n141 ) : ( 10'd640 ) ;
assign n143 =  ( n34 ) ? ( LB2D_shift_y ) : ( LB2D_shift_y ) ;
assign n144 =  ( n27 ) ? ( LB2D_shift_y ) : ( n143 ) ;
assign n145 =  ( n22 ) ? ( n142 ) : ( n144 ) ;
assign n146 =  ( n13 ) ? ( LB2D_shift_y ) : ( n145 ) ;
assign n147 =  ( n4 ) ? ( LB2D_shift_y ) : ( n146 ) ;
assign n148 =  ( stencil_stream_full ) == ( 1'd1 )  ;
assign n149 =  ( n148 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_0 ) ;
//assign n150 = gb_fun(n149) ;
gb_fun gb_fun_U (
        .a (n149),
        .b (n150)
        );

assign n151 =  ( n34 ) ? ( arg_0_TDATA ) : ( arg_0_TDATA ) ;
assign n152 =  ( n27 ) ? ( arg_0_TDATA ) : ( n151 ) ;
assign n153 =  ( n22 ) ? ( arg_0_TDATA ) : ( n152 ) ;
assign n154 =  ( n13 ) ? ( n150 ) : ( n153 ) ;
assign n155 =  ( n4 ) ? ( arg_0_TDATA ) : ( n154 ) ;
assign n156 =  ( gb_pp_it_8 ) == ( 1'd1 )  ;
assign n157 =  ( n156 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n158 =  ( n34 ) ? ( arg_0_TVALID ) : ( arg_0_TVALID ) ;
assign n159 =  ( n27 ) ? ( arg_0_TVALID ) : ( n158 ) ;
assign n160 =  ( n22 ) ? ( arg_0_TVALID ) : ( n159 ) ;
assign n161 =  ( n13 ) ? ( n157 ) : ( n160 ) ;
assign n162 =  ( n4 ) ? ( 1'd0 ) : ( n161 ) ;
assign n163 =  ( 19'd316224 ) - ( 19'd1 )  ;
assign n164 =  ( LB1D_p_cnt ) == ( n163 )  ;
assign n165 =  ( n164 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n166 =  ( n34 ) ? ( n165 ) : ( arg_1_TREADY ) ;
assign n167 =  ( n32 ) ? ( 1'd1 ) : ( n166 ) ;
assign n168 =  ( n27 ) ? ( arg_1_TREADY ) : ( n167 ) ;
assign n169 =  ( n22 ) ? ( arg_1_TREADY ) : ( n168 ) ;
assign n170 =  ( n13 ) ? ( arg_1_TREADY ) : ( n169 ) ;
assign n171 =  ( n4 ) ? ( arg_1_TREADY ) : ( n170 ) ;
assign n172 =  ( gb_p_cnt ) + ( 19'd1 )  ;
assign n173 =  ( n172 ) == ( 19'd307200 )  ;
assign n174 =  ( n173 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n175 =  ( n34 ) ? ( gb_exit_it_1 ) : ( gb_exit_it_1 ) ;
assign n176 =  ( n27 ) ? ( gb_exit_it_1 ) : ( n175 ) ;
assign n177 =  ( n22 ) ? ( gb_exit_it_1 ) : ( n176 ) ;
assign n178 =  ( n13 ) ? ( n174 ) : ( n177 ) ;
assign n179 =  ( n4 ) ? ( gb_exit_it_1 ) : ( n178 ) ;
assign n180 =  ( n34 ) ? ( gb_exit_it_2 ) : ( gb_exit_it_2 ) ;
assign n181 =  ( n27 ) ? ( gb_exit_it_2 ) : ( n180 ) ;
assign n182 =  ( n22 ) ? ( gb_exit_it_2 ) : ( n181 ) ;
assign n183 =  ( n13 ) ? ( gb_exit_it_1 ) : ( n182 ) ;
assign n184 =  ( n4 ) ? ( gb_exit_it_2 ) : ( n183 ) ;
assign n185 =  ( n34 ) ? ( gb_exit_it_3 ) : ( gb_exit_it_3 ) ;
assign n186 =  ( n27 ) ? ( gb_exit_it_3 ) : ( n185 ) ;
assign n187 =  ( n22 ) ? ( gb_exit_it_3 ) : ( n186 ) ;
assign n188 =  ( n13 ) ? ( gb_exit_it_2 ) : ( n187 ) ;
assign n189 =  ( n4 ) ? ( gb_exit_it_3 ) : ( n188 ) ;
assign n190 =  ( n34 ) ? ( gb_exit_it_4 ) : ( gb_exit_it_4 ) ;
assign n191 =  ( n27 ) ? ( gb_exit_it_4 ) : ( n190 ) ;
assign n192 =  ( n22 ) ? ( gb_exit_it_4 ) : ( n191 ) ;
assign n193 =  ( n13 ) ? ( gb_exit_it_3 ) : ( n192 ) ;
assign n194 =  ( n4 ) ? ( gb_exit_it_4 ) : ( n193 ) ;
assign n195 =  ( n34 ) ? ( gb_exit_it_5 ) : ( gb_exit_it_5 ) ;
assign n196 =  ( n27 ) ? ( gb_exit_it_5 ) : ( n195 ) ;
assign n197 =  ( n22 ) ? ( gb_exit_it_5 ) : ( n196 ) ;
assign n198 =  ( n13 ) ? ( gb_exit_it_4 ) : ( n197 ) ;
assign n199 =  ( n4 ) ? ( gb_exit_it_5 ) : ( n198 ) ;
assign n200 =  ( n34 ) ? ( gb_exit_it_6 ) : ( gb_exit_it_6 ) ;
assign n201 =  ( n27 ) ? ( gb_exit_it_6 ) : ( n200 ) ;
assign n202 =  ( n22 ) ? ( gb_exit_it_6 ) : ( n201 ) ;
assign n203 =  ( n13 ) ? ( gb_exit_it_5 ) : ( n202 ) ;
assign n204 =  ( n4 ) ? ( gb_exit_it_6 ) : ( n203 ) ;
assign n205 =  ( n34 ) ? ( gb_exit_it_7 ) : ( gb_exit_it_7 ) ;
assign n206 =  ( n27 ) ? ( gb_exit_it_7 ) : ( n205 ) ;
assign n207 =  ( n22 ) ? ( gb_exit_it_7 ) : ( n206 ) ;
assign n208 =  ( n13 ) ? ( gb_exit_it_6 ) : ( n207 ) ;
assign n209 =  ( n4 ) ? ( gb_exit_it_7 ) : ( n208 ) ;
assign n210 =  ( n34 ) ? ( gb_exit_it_8 ) : ( gb_exit_it_8 ) ;
assign n211 =  ( n27 ) ? ( gb_exit_it_8 ) : ( n210 ) ;
assign n212 =  ( n22 ) ? ( gb_exit_it_8 ) : ( n211 ) ;
assign n213 =  ( n13 ) ? ( gb_exit_it_7 ) : ( n212 ) ;
assign n214 =  ( n4 ) ? ( gb_exit_it_8 ) : ( n213 ) ;
assign n215 =  ( gb_p_cnt ) < ( 19'd307200 )  ;
assign n216 =  ( n215 ) ? ( n172 ) : ( 19'd307200 ) ;
assign n217 =  ( n34 ) ? ( gb_p_cnt ) : ( gb_p_cnt ) ;
assign n218 =  ( n27 ) ? ( gb_p_cnt ) : ( n217 ) ;
assign n219 =  ( n22 ) ? ( gb_p_cnt ) : ( n218 ) ;
assign n220 =  ( n13 ) ? ( n216 ) : ( n219 ) ;
assign n221 =  ( n4 ) ? ( gb_p_cnt ) : ( n220 ) ;
assign n222 =  ( n34 ) ? ( gb_pp_it_1 ) : ( gb_pp_it_1 ) ;
assign n223 =  ( n27 ) ? ( gb_pp_it_1 ) : ( n222 ) ;
assign n224 =  ( n22 ) ? ( gb_pp_it_1 ) : ( n223 ) ;
assign n225 =  ( n13 ) ? ( 1'd1 ) : ( n224 ) ;
assign n226 =  ( n4 ) ? ( gb_pp_it_1 ) : ( n225 ) ;
assign n227 =  ( n34 ) ? ( gb_pp_it_2 ) : ( gb_pp_it_2 ) ;
assign n228 =  ( n27 ) ? ( gb_pp_it_2 ) : ( n227 ) ;
assign n229 =  ( n22 ) ? ( gb_pp_it_2 ) : ( n228 ) ;
assign n230 =  ( n13 ) ? ( gb_pp_it_1 ) : ( n229 ) ;
assign n231 =  ( n4 ) ? ( gb_pp_it_2 ) : ( n230 ) ;
assign n232 =  ( n34 ) ? ( gb_pp_it_3 ) : ( gb_pp_it_3 ) ;
assign n233 =  ( n27 ) ? ( gb_pp_it_3 ) : ( n232 ) ;
assign n234 =  ( n22 ) ? ( gb_pp_it_3 ) : ( n233 ) ;
assign n235 =  ( n13 ) ? ( gb_pp_it_2 ) : ( n234 ) ;
assign n236 =  ( n4 ) ? ( gb_pp_it_3 ) : ( n235 ) ;
assign n237 =  ( n34 ) ? ( gb_pp_it_4 ) : ( gb_pp_it_4 ) ;
assign n238 =  ( n27 ) ? ( gb_pp_it_4 ) : ( n237 ) ;
assign n239 =  ( n22 ) ? ( gb_pp_it_4 ) : ( n238 ) ;
assign n240 =  ( n13 ) ? ( gb_pp_it_3 ) : ( n239 ) ;
assign n241 =  ( n4 ) ? ( gb_pp_it_4 ) : ( n240 ) ;
assign n242 =  ( n34 ) ? ( gb_pp_it_5 ) : ( gb_pp_it_5 ) ;
assign n243 =  ( n27 ) ? ( gb_pp_it_5 ) : ( n242 ) ;
assign n244 =  ( n22 ) ? ( gb_pp_it_5 ) : ( n243 ) ;
assign n245 =  ( n13 ) ? ( gb_pp_it_4 ) : ( n244 ) ;
assign n246 =  ( n4 ) ? ( gb_pp_it_5 ) : ( n245 ) ;
assign n247 =  ( n34 ) ? ( gb_pp_it_6 ) : ( gb_pp_it_6 ) ;
assign n248 =  ( n27 ) ? ( gb_pp_it_6 ) : ( n247 ) ;
assign n249 =  ( n22 ) ? ( gb_pp_it_6 ) : ( n248 ) ;
assign n250 =  ( n13 ) ? ( gb_pp_it_5 ) : ( n249 ) ;
assign n251 =  ( n4 ) ? ( gb_pp_it_6 ) : ( n250 ) ;
assign n252 =  ( n34 ) ? ( gb_pp_it_7 ) : ( gb_pp_it_7 ) ;
assign n253 =  ( n27 ) ? ( gb_pp_it_7 ) : ( n252 ) ;
assign n254 =  ( n22 ) ? ( gb_pp_it_7 ) : ( n253 ) ;
assign n255 =  ( n13 ) ? ( gb_pp_it_6 ) : ( n254 ) ;
assign n256 =  ( n4 ) ? ( gb_pp_it_7 ) : ( n255 ) ;
assign n257 =  ( n34 ) ? ( gb_pp_it_8 ) : ( gb_pp_it_8 ) ;
assign n258 =  ( n27 ) ? ( gb_pp_it_8 ) : ( n257 ) ;
assign n259 =  ( n22 ) ? ( gb_pp_it_8 ) : ( n258 ) ;
assign n260 =  ( n13 ) ? ( gb_pp_it_7 ) : ( n259 ) ;
assign n261 =  ( n4 ) ? ( gb_pp_it_8 ) : ( n260 ) ;
assign n262 =  ( n34 ) ? ( gb_pp_it_9 ) : ( gb_pp_it_9 ) ;
assign n263 =  ( n27 ) ? ( gb_pp_it_9 ) : ( n262 ) ;
assign n264 =  ( n22 ) ? ( gb_pp_it_9 ) : ( n263 ) ;
assign n265 =  ( n13 ) ? ( gb_pp_it_8 ) : ( n264 ) ;
assign n266 =  ( n4 ) ? ( gb_pp_it_9 ) : ( n265 ) ;
assign n267 =  ( n34 ) ? ( LB1D_uIn ) : ( in_stream_buff_0 ) ;
assign n268 =  ( n27 ) ? ( in_stream_buff_0 ) : ( n267 ) ;
assign n269 =  ( n22 ) ? ( in_stream_buff_0 ) : ( n268 ) ;
assign n270 =  ( n13 ) ? ( in_stream_buff_0 ) : ( n269 ) ;
assign n271 =  ( n4 ) ? ( in_stream_buff_0 ) : ( n270 ) ;
assign n272 =  ( n34 ) ? ( in_stream_buff_0 ) : ( in_stream_buff_1 ) ;
assign n273 =  ( n27 ) ? ( in_stream_buff_1 ) : ( n272 ) ;
assign n274 =  ( n22 ) ? ( in_stream_buff_1 ) : ( n273 ) ;
assign n275 =  ( n13 ) ? ( in_stream_buff_1 ) : ( n274 ) ;
assign n276 =  ( n4 ) ? ( in_stream_buff_1 ) : ( n275 ) ;
assign n277 =  ( in_stream_full ) == ( 1'd1 )  ;
assign n278 =  ( n277 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n279 =  ( n34 ) ? ( 1'd0 ) : ( in_stream_empty ) ;
assign n280 =  ( n27 ) ? ( n278 ) : ( n279 ) ;
assign n281 =  ( n22 ) ? ( in_stream_empty ) : ( n280 ) ;
assign n282 =  ( n13 ) ? ( in_stream_empty ) : ( n281 ) ;
assign n283 =  ( n4 ) ? ( in_stream_empty ) : ( n282 ) ;
assign n284 =  ( in_stream_empty ) == ( 1'd1 )  ;
assign n285 =  ( n284 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n286 =  ( n34 ) ? ( n285 ) : ( in_stream_full ) ;
assign n287 =  ( n27 ) ? ( 1'd0 ) : ( n286 ) ;
assign n288 =  ( n22 ) ? ( in_stream_full ) : ( n287 ) ;
assign n289 =  ( n13 ) ? ( in_stream_full ) : ( n288 ) ;
assign n290 =  ( n4 ) ? ( in_stream_full ) : ( n289 ) ;
assign n291 =  ( n277 ) ? ( in_stream_buff_1 ) : ( in_stream_buff_0 ) ;
assign n292 =  ( LB2D_proc_w ) == ( 64'd0 )  ;
assign n293 =  ( LB2D_proc_x ) - ( 9'd1 )  ;
assign n294 =  (  LB2D_proc_7 [ n293 ] )  ;
assign n295 =  ( LB2D_proc_w ) == ( 64'd1 )  ;
assign n296 =  (  LB2D_proc_0 [ n293 ] )  ;
assign n297 =  ( LB2D_proc_w ) == ( 64'd2 )  ;
assign n298 =  (  LB2D_proc_1 [ n293 ] )  ;
assign n299 =  ( LB2D_proc_w ) == ( 64'd3 )  ;
assign n300 =  (  LB2D_proc_2 [ n293 ] )  ;
assign n301 =  ( LB2D_proc_w ) == ( 64'd4 )  ;
assign n302 =  (  LB2D_proc_3 [ n293 ] )  ;
assign n303 =  ( LB2D_proc_w ) == ( 64'd5 )  ;
assign n304 =  (  LB2D_proc_4 [ n293 ] )  ;
assign n305 =  ( LB2D_proc_w ) == ( 64'd6 )  ;
assign n306 =  (  LB2D_proc_5 [ n293 ] )  ;
assign n307 =  (  LB2D_proc_6 [ n293 ] )  ;
assign n308 =  ( n305 ) ? ( n306 ) : ( n307 ) ;
assign n309 =  ( n303 ) ? ( n304 ) : ( n308 ) ;
assign n310 =  ( n301 ) ? ( n302 ) : ( n309 ) ;
assign n311 =  ( n299 ) ? ( n300 ) : ( n310 ) ;
assign n312 =  ( n297 ) ? ( n298 ) : ( n311 ) ;
assign n313 =  ( n295 ) ? ( n296 ) : ( n312 ) ;
assign n314 =  ( n292 ) ? ( n294 ) : ( n313 ) ;
assign n315 =  ( n305 ) ? ( n304 ) : ( n306 ) ;
assign n316 =  ( n303 ) ? ( n302 ) : ( n315 ) ;
assign n317 =  ( n301 ) ? ( n300 ) : ( n316 ) ;
assign n318 =  ( n299 ) ? ( n298 ) : ( n317 ) ;
assign n319 =  ( n297 ) ? ( n296 ) : ( n318 ) ;
assign n320 =  ( n295 ) ? ( n294 ) : ( n319 ) ;
assign n321 =  ( n292 ) ? ( n307 ) : ( n320 ) ;
assign n322 =  ( n305 ) ? ( n302 ) : ( n304 ) ;
assign n323 =  ( n303 ) ? ( n300 ) : ( n322 ) ;
assign n324 =  ( n301 ) ? ( n298 ) : ( n323 ) ;
assign n325 =  ( n299 ) ? ( n296 ) : ( n324 ) ;
assign n326 =  ( n297 ) ? ( n294 ) : ( n325 ) ;
assign n327 =  ( n295 ) ? ( n307 ) : ( n326 ) ;
assign n328 =  ( n292 ) ? ( n306 ) : ( n327 ) ;
assign n329 =  ( n305 ) ? ( n300 ) : ( n302 ) ;
assign n330 =  ( n303 ) ? ( n298 ) : ( n329 ) ;
assign n331 =  ( n301 ) ? ( n296 ) : ( n330 ) ;
assign n332 =  ( n299 ) ? ( n294 ) : ( n331 ) ;
assign n333 =  ( n297 ) ? ( n307 ) : ( n332 ) ;
assign n334 =  ( n295 ) ? ( n306 ) : ( n333 ) ;
assign n335 =  ( n292 ) ? ( n304 ) : ( n334 ) ;
assign n336 =  ( n305 ) ? ( n298 ) : ( n300 ) ;
assign n337 =  ( n303 ) ? ( n296 ) : ( n336 ) ;
assign n338 =  ( n301 ) ? ( n294 ) : ( n337 ) ;
assign n339 =  ( n299 ) ? ( n307 ) : ( n338 ) ;
assign n340 =  ( n297 ) ? ( n306 ) : ( n339 ) ;
assign n341 =  ( n295 ) ? ( n304 ) : ( n340 ) ;
assign n342 =  ( n292 ) ? ( n302 ) : ( n341 ) ;
assign n343 =  ( n305 ) ? ( n296 ) : ( n298 ) ;
assign n344 =  ( n303 ) ? ( n294 ) : ( n343 ) ;
assign n345 =  ( n301 ) ? ( n307 ) : ( n344 ) ;
assign n346 =  ( n299 ) ? ( n306 ) : ( n345 ) ;
assign n347 =  ( n297 ) ? ( n304 ) : ( n346 ) ;
assign n348 =  ( n295 ) ? ( n302 ) : ( n347 ) ;
assign n349 =  ( n292 ) ? ( n300 ) : ( n348 ) ;
assign n350 =  ( n305 ) ? ( n294 ) : ( n296 ) ;
assign n351 =  ( n303 ) ? ( n307 ) : ( n350 ) ;
assign n352 =  ( n301 ) ? ( n306 ) : ( n351 ) ;
assign n353 =  ( n299 ) ? ( n304 ) : ( n352 ) ;
assign n354 =  ( n297 ) ? ( n302 ) : ( n353 ) ;
assign n355 =  ( n295 ) ? ( n300 ) : ( n354 ) ;
assign n356 =  ( n292 ) ? ( n298 ) : ( n355 ) ;
assign n357 =  ( n305 ) ? ( n307 ) : ( n294 ) ;
assign n358 =  ( n303 ) ? ( n306 ) : ( n357 ) ;
assign n359 =  ( n301 ) ? ( n304 ) : ( n358 ) ;
assign n360 =  ( n299 ) ? ( n302 ) : ( n359 ) ;
assign n361 =  ( n297 ) ? ( n300 ) : ( n360 ) ;
assign n362 =  ( n295 ) ? ( n298 ) : ( n361 ) ;
assign n363 =  ( n292 ) ? ( n296 ) : ( n362 ) ;
assign n364 =  { ( n356 ) , ( n363 ) }  ;
assign n365 =  { ( n349 ) , ( n364 ) }  ;
assign n366 =  { ( n342 ) , ( n365 ) }  ;
assign n367 =  { ( n335 ) , ( n366 ) }  ;
assign n368 =  { ( n328 ) , ( n367 ) }  ;
assign n369 =  { ( n321 ) , ( n368 ) }  ;
assign n370 =  { ( n314 ) , ( n369 ) }  ;
assign n371 =  { ( n291 ) , ( n370 ) }  ;
assign n372 =  ( n25 ) ? ( slice_stream_buff_0 ) : ( n371 ) ;
assign n373 =  ( n34 ) ? ( slice_stream_buff_0 ) : ( slice_stream_buff_0 ) ;
assign n374 =  ( n27 ) ? ( n372 ) : ( n373 ) ;
assign n375 =  ( n22 ) ? ( slice_stream_buff_0 ) : ( n374 ) ;
assign n376 =  ( n13 ) ? ( slice_stream_buff_0 ) : ( n375 ) ;
assign n377 =  ( n4 ) ? ( slice_stream_buff_0 ) : ( n376 ) ;
assign n378 =  ( n25 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n379 =  ( n34 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_1 ) ;
assign n380 =  ( n27 ) ? ( n378 ) : ( n379 ) ;
assign n381 =  ( n22 ) ? ( slice_stream_buff_1 ) : ( n380 ) ;
assign n382 =  ( n13 ) ? ( slice_stream_buff_1 ) : ( n381 ) ;
assign n383 =  ( n4 ) ? ( slice_stream_buff_1 ) : ( n382 ) ;
assign n384 =  ( n125 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n385 =  ( n25 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n386 =  ( n34 ) ? ( slice_stream_empty ) : ( slice_stream_empty ) ;
assign n387 =  ( n27 ) ? ( n385 ) : ( n386 ) ;
assign n388 =  ( n22 ) ? ( n384 ) : ( n387 ) ;
assign n389 =  ( n13 ) ? ( slice_stream_empty ) : ( n388 ) ;
assign n390 =  ( n4 ) ? ( slice_stream_empty ) : ( n389 ) ;
assign n391 =  ( slice_stream_empty ) == ( 1'd1 )  ;
assign n392 =  ( n391 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n393 =  ( n25 ) ? ( 1'd0 ) : ( n392 ) ;
assign n394 =  ( n34 ) ? ( slice_stream_full ) : ( slice_stream_full ) ;
assign n395 =  ( n27 ) ? ( n393 ) : ( n394 ) ;
assign n396 =  ( n22 ) ? ( 1'd0 ) : ( n395 ) ;
assign n397 =  ( n13 ) ? ( slice_stream_full ) : ( n396 ) ;
assign n398 =  ( n4 ) ? ( slice_stream_full ) : ( n397 ) ;
assign n399 =  ( LB2D_shift_x ) >= ( 9'd8 )  ;
assign n400 =  ( LB2D_shift_x ) == ( 9'd0 )  ;
assign n401 =  ( n399 ) | ( n400 )  ;
assign n402 = n126[71:64] ;
assign n403 = LB2D_shift_7[71:64] ;
assign n404 = LB2D_shift_6[71:64] ;
assign n405 = LB2D_shift_5[71:64] ;
assign n406 = LB2D_shift_4[71:64] ;
assign n407 = LB2D_shift_3[71:64] ;
assign n408 = LB2D_shift_2[71:64] ;
assign n409 = LB2D_shift_1[71:64] ;
assign n410 = LB2D_shift_0[71:64] ;
assign n411 =  { ( n409 ) , ( n410 ) }  ;
assign n412 =  { ( n408 ) , ( n411 ) }  ;
assign n413 =  { ( n407 ) , ( n412 ) }  ;
assign n414 =  { ( n406 ) , ( n413 ) }  ;
assign n415 =  { ( n405 ) , ( n414 ) }  ;
assign n416 =  { ( n404 ) , ( n415 ) }  ;
assign n417 =  { ( n403 ) , ( n416 ) }  ;
assign n418 =  { ( n402 ) , ( n417 ) }  ;
assign n419 = n126[63:56] ;
assign n420 = LB2D_shift_7[63:56] ;
assign n421 = LB2D_shift_6[63:56] ;
assign n422 = LB2D_shift_5[63:56] ;
assign n423 = LB2D_shift_4[63:56] ;
assign n424 = LB2D_shift_3[63:56] ;
assign n425 = LB2D_shift_2[63:56] ;
assign n426 = LB2D_shift_1[63:56] ;
assign n427 = LB2D_shift_0[63:56] ;
assign n428 =  { ( n426 ) , ( n427 ) }  ;
assign n429 =  { ( n425 ) , ( n428 ) }  ;
assign n430 =  { ( n424 ) , ( n429 ) }  ;
assign n431 =  { ( n423 ) , ( n430 ) }  ;
assign n432 =  { ( n422 ) , ( n431 ) }  ;
assign n433 =  { ( n421 ) , ( n432 ) }  ;
assign n434 =  { ( n420 ) , ( n433 ) }  ;
assign n435 =  { ( n419 ) , ( n434 ) }  ;
assign n436 = n126[55:48] ;
assign n437 = LB2D_shift_7[55:48] ;
assign n438 = LB2D_shift_6[55:48] ;
assign n439 = LB2D_shift_5[55:48] ;
assign n440 = LB2D_shift_4[55:48] ;
assign n441 = LB2D_shift_3[55:48] ;
assign n442 = LB2D_shift_2[55:48] ;
assign n443 = LB2D_shift_1[55:48] ;
assign n444 = LB2D_shift_0[55:48] ;
assign n445 =  { ( n443 ) , ( n444 ) }  ;
assign n446 =  { ( n442 ) , ( n445 ) }  ;
assign n447 =  { ( n441 ) , ( n446 ) }  ;
assign n448 =  { ( n440 ) , ( n447 ) }  ;
assign n449 =  { ( n439 ) , ( n448 ) }  ;
assign n450 =  { ( n438 ) , ( n449 ) }  ;
assign n451 =  { ( n437 ) , ( n450 ) }  ;
assign n452 =  { ( n436 ) , ( n451 ) }  ;
assign n453 = n126[47:40] ;
assign n454 = LB2D_shift_7[47:40] ;
assign n455 = LB2D_shift_6[47:40] ;
assign n456 = LB2D_shift_5[47:40] ;
assign n457 = LB2D_shift_4[47:40] ;
assign n458 = LB2D_shift_3[47:40] ;
assign n459 = LB2D_shift_2[47:40] ;
assign n460 = LB2D_shift_1[47:40] ;
assign n461 = LB2D_shift_0[47:40] ;
assign n462 =  { ( n460 ) , ( n461 ) }  ;
assign n463 =  { ( n459 ) , ( n462 ) }  ;
assign n464 =  { ( n458 ) , ( n463 ) }  ;
assign n465 =  { ( n457 ) , ( n464 ) }  ;
assign n466 =  { ( n456 ) , ( n465 ) }  ;
assign n467 =  { ( n455 ) , ( n466 ) }  ;
assign n468 =  { ( n454 ) , ( n467 ) }  ;
assign n469 =  { ( n453 ) , ( n468 ) }  ;
assign n470 = n126[39:32] ;
assign n471 = LB2D_shift_7[39:32] ;
assign n472 = LB2D_shift_6[39:32] ;
assign n473 = LB2D_shift_5[39:32] ;
assign n474 = LB2D_shift_4[39:32] ;
assign n475 = LB2D_shift_3[39:32] ;
assign n476 = LB2D_shift_2[39:32] ;
assign n477 = LB2D_shift_1[39:32] ;
assign n478 = LB2D_shift_0[39:32] ;
assign n479 =  { ( n477 ) , ( n478 ) }  ;
assign n480 =  { ( n476 ) , ( n479 ) }  ;
assign n481 =  { ( n475 ) , ( n480 ) }  ;
assign n482 =  { ( n474 ) , ( n481 ) }  ;
assign n483 =  { ( n473 ) , ( n482 ) }  ;
assign n484 =  { ( n472 ) , ( n483 ) }  ;
assign n485 =  { ( n471 ) , ( n484 ) }  ;
assign n486 =  { ( n470 ) , ( n485 ) }  ;
assign n487 = n126[31:24] ;
assign n488 = LB2D_shift_7[31:24] ;
assign n489 = LB2D_shift_6[31:24] ;
assign n490 = LB2D_shift_5[31:24] ;
assign n491 = LB2D_shift_4[31:24] ;
assign n492 = LB2D_shift_3[31:24] ;
assign n493 = LB2D_shift_2[31:24] ;
assign n494 = LB2D_shift_1[31:24] ;
assign n495 = LB2D_shift_0[31:24] ;
assign n496 =  { ( n494 ) , ( n495 ) }  ;
assign n497 =  { ( n493 ) , ( n496 ) }  ;
assign n498 =  { ( n492 ) , ( n497 ) }  ;
assign n499 =  { ( n491 ) , ( n498 ) }  ;
assign n500 =  { ( n490 ) , ( n499 ) }  ;
assign n501 =  { ( n489 ) , ( n500 ) }  ;
assign n502 =  { ( n488 ) , ( n501 ) }  ;
assign n503 =  { ( n487 ) , ( n502 ) }  ;
assign n504 = n126[23:16] ;
assign n505 = LB2D_shift_7[23:16] ;
assign n506 = LB2D_shift_6[23:16] ;
assign n507 = LB2D_shift_5[23:16] ;
assign n508 = LB2D_shift_4[23:16] ;
assign n509 = LB2D_shift_3[23:16] ;
assign n510 = LB2D_shift_2[23:16] ;
assign n511 = LB2D_shift_1[23:16] ;
assign n512 = LB2D_shift_0[23:16] ;
assign n513 =  { ( n511 ) , ( n512 ) }  ;
assign n514 =  { ( n510 ) , ( n513 ) }  ;
assign n515 =  { ( n509 ) , ( n514 ) }  ;
assign n516 =  { ( n508 ) , ( n515 ) }  ;
assign n517 =  { ( n507 ) , ( n516 ) }  ;
assign n518 =  { ( n506 ) , ( n517 ) }  ;
assign n519 =  { ( n505 ) , ( n518 ) }  ;
assign n520 =  { ( n504 ) , ( n519 ) }  ;
assign n521 = n126[15:8] ;
assign n522 = LB2D_shift_7[15:8] ;
assign n523 = LB2D_shift_6[15:8] ;
assign n524 = LB2D_shift_5[15:8] ;
assign n525 = LB2D_shift_4[15:8] ;
assign n526 = LB2D_shift_3[15:8] ;
assign n527 = LB2D_shift_2[15:8] ;
assign n528 = LB2D_shift_1[15:8] ;
assign n529 = LB2D_shift_0[15:8] ;
assign n530 =  { ( n528 ) , ( n529 ) }  ;
assign n531 =  { ( n527 ) , ( n530 ) }  ;
assign n532 =  { ( n526 ) , ( n531 ) }  ;
assign n533 =  { ( n525 ) , ( n532 ) }  ;
assign n534 =  { ( n524 ) , ( n533 ) }  ;
assign n535 =  { ( n523 ) , ( n534 ) }  ;
assign n536 =  { ( n522 ) , ( n535 ) }  ;
assign n537 =  { ( n521 ) , ( n536 ) }  ;
assign n538 = n126[7:0] ;
assign n539 = LB2D_shift_7[7:0] ;
assign n540 = LB2D_shift_6[7:0] ;
assign n541 = LB2D_shift_5[7:0] ;
assign n542 = LB2D_shift_4[7:0] ;
assign n543 = LB2D_shift_3[7:0] ;
assign n544 = LB2D_shift_2[7:0] ;
assign n545 = LB2D_shift_1[7:0] ;
assign n546 = LB2D_shift_0[7:0] ;
assign n547 =  { ( n545 ) , ( n546 ) }  ;
assign n548 =  { ( n544 ) , ( n547 ) }  ;
assign n549 =  { ( n543 ) , ( n548 ) }  ;
assign n550 =  { ( n542 ) , ( n549 ) }  ;
assign n551 =  { ( n541 ) , ( n550 ) }  ;
assign n552 =  { ( n540 ) , ( n551 ) }  ;
assign n553 =  { ( n539 ) , ( n552 ) }  ;
assign n554 =  { ( n538 ) , ( n553 ) }  ;
assign n555 =  { ( n537 ) , ( n554 ) }  ;
assign n556 =  { ( n520 ) , ( n555 ) }  ;
assign n557 =  { ( n503 ) , ( n556 ) }  ;
assign n558 =  { ( n486 ) , ( n557 ) }  ;
assign n559 =  { ( n469 ) , ( n558 ) }  ;
assign n560 =  { ( n452 ) , ( n559 ) }  ;
assign n561 =  { ( n435 ) , ( n560 ) }  ;
assign n562 =  { ( n418 ) , ( n561 ) }  ;
assign n563 =  ( n401 ) ? ( n562 ) : ( stencil_stream_buff_0 ) ;
assign n564 =  ( n34 ) ? ( stencil_stream_buff_0 ) : ( stencil_stream_buff_0 ) ;
assign n565 =  ( n27 ) ? ( stencil_stream_buff_0 ) : ( n564 ) ;
assign n566 =  ( n22 ) ? ( n563 ) : ( n565 ) ;
assign n567 =  ( n13 ) ? ( stencil_stream_buff_0 ) : ( n566 ) ;
assign n568 =  ( n4 ) ? ( stencil_stream_buff_0 ) : ( n567 ) ;
assign n569 =  ( n34 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_1 ) ;
assign n570 =  ( n27 ) ? ( stencil_stream_buff_1 ) : ( n569 ) ;
assign n571 =  ( n22 ) ? ( stencil_stream_buff_0 ) : ( n570 ) ;
assign n572 =  ( n13 ) ? ( stencil_stream_buff_1 ) : ( n571 ) ;
assign n573 =  ( n4 ) ? ( stencil_stream_buff_1 ) : ( n572 ) ;
assign n574 =  ( n148 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n575 = ~ ( n401 ) ;
assign n576 =  ( n575 ) ? ( stencil_stream_empty ) : ( 1'd0 ) ;
assign n577 =  ( n34 ) ? ( stencil_stream_empty ) : ( stencil_stream_empty ) ;
assign n578 =  ( n27 ) ? ( stencil_stream_empty ) : ( n577 ) ;
assign n579 =  ( n22 ) ? ( n576 ) : ( n578 ) ;
assign n580 =  ( n13 ) ? ( n574 ) : ( n579 ) ;
assign n581 =  ( n4 ) ? ( stencil_stream_empty ) : ( n580 ) ;
assign n582 =  ( n9 ) ? ( 1'd0 ) : ( 1'd0 ) ;
assign n583 =  ( stencil_stream_empty ) == ( 1'd1 )  ;
assign n584 =  ( n583 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n585 =  ( n575 ) ? ( stencil_stream_full ) : ( n584 ) ;
assign n586 =  ( n34 ) ? ( stencil_stream_full ) : ( stencil_stream_full ) ;
assign n587 =  ( n27 ) ? ( stencil_stream_full ) : ( n586 ) ;
assign n588 =  ( n22 ) ? ( n585 ) : ( n587 ) ;
assign n589 =  ( n13 ) ? ( n582 ) : ( n588 ) ;
assign n590 =  ( n4 ) ? ( stencil_stream_full ) : ( n589 ) ;
assign n591 = ~ ( n4 ) ;
assign n592 = ~ ( n13 ) ;
assign n593 =  ( n591 ) & ( n592 )  ;
assign n594 = ~ ( n22 ) ;
assign n595 =  ( n593 ) & ( n594 )  ;
assign n596 = ~ ( n27 ) ;
assign n597 =  ( n595 ) & ( n596 )  ;
assign n598 = ~ ( n34 ) ;
assign n599 =  ( n597 ) & ( n598 )  ;
assign n600 =  ( n597 ) & ( n34 )  ;
assign n601 =  ( n595 ) & ( n27 )  ;
assign n602 = ~ ( n292 ) ;
assign n603 =  ( n601 ) & ( n602 )  ;
assign n604 =  ( n601 ) & ( n292 )  ;
assign n605 =  ( n593 ) & ( n22 )  ;
assign n606 =  ( n591 ) & ( n13 )  ;
assign LB2D_proc_0_addr0 = n604 ? (n293) : (0);
assign LB2D_proc_0_data0 = n604 ? (n291) : (LB2D_proc_0[0]);
assign n607 = ~ ( n295 ) ;
assign n608 =  ( n601 ) & ( n607 )  ;
assign n609 =  ( n601 ) & ( n295 )  ;
assign LB2D_proc_1_addr0 = n609 ? (n293) : (0);
assign LB2D_proc_1_data0 = n609 ? (n291) : (LB2D_proc_1[0]);
assign n610 = ~ ( n297 ) ;
assign n611 =  ( n601 ) & ( n610 )  ;
assign n612 =  ( n601 ) & ( n297 )  ;
assign LB2D_proc_2_addr0 = n612 ? (n293) : (0);
assign LB2D_proc_2_data0 = n612 ? (n291) : (LB2D_proc_2[0]);
assign n613 = ~ ( n299 ) ;
assign n614 =  ( n601 ) & ( n613 )  ;
assign n615 =  ( n601 ) & ( n299 )  ;
assign LB2D_proc_3_addr0 = n615 ? (n293) : (0);
assign LB2D_proc_3_data0 = n615 ? (n291) : (LB2D_proc_3[0]);
assign n616 = ~ ( n301 ) ;
assign n617 =  ( n601 ) & ( n616 )  ;
assign n618 =  ( n601 ) & ( n301 )  ;
assign LB2D_proc_4_addr0 = n618 ? (n293) : (0);
assign LB2D_proc_4_data0 = n618 ? (n291) : (LB2D_proc_4[0]);
assign n619 = ~ ( n303 ) ;
assign n620 =  ( n601 ) & ( n619 )  ;
assign n621 =  ( n601 ) & ( n303 )  ;
assign LB2D_proc_5_addr0 = n621 ? (n293) : (0);
assign LB2D_proc_5_data0 = n621 ? (n291) : (LB2D_proc_5[0]);
assign n622 = ~ ( n305 ) ;
assign n623 =  ( n601 ) & ( n622 )  ;
assign n624 =  ( n601 ) & ( n305 )  ;
assign LB2D_proc_6_addr0 = n624 ? (n293) : (0);
assign LB2D_proc_6_data0 = n624 ? (n291) : (LB2D_proc_6[0]);
assign n625 = ~ ( n65 ) ;
assign n626 =  ( n601 ) & ( n625 )  ;
assign n627 =  ( n601 ) & ( n65 )  ;
assign LB2D_proc_7_addr0 = n627 ? (n293) : (0);
assign LB2D_proc_7_data0 = n627 ? (n291) : (LB2D_proc_7[0]);
/*
function [7:0] gb_fun ;
input [647:0] arg0;
    begin
//TODO: Add the specific function HERE.    end
endfunction
*/

always @(posedge clk) begin
   if(rst) begin
       LB1D_buff <= LB1D_buff;
       LB1D_in <= LB1D_in;
       LB1D_it_1 <= LB1D_it_1;
       LB1D_p_cnt <= LB1D_p_cnt;
       LB1D_uIn <= LB1D_uIn;
       LB2D_proc_w <= LB2D_proc_w;
       LB2D_proc_x <= LB2D_proc_x;
       LB2D_proc_y <= LB2D_proc_y;
       LB2D_shift_0 <= LB2D_shift_0;
       LB2D_shift_1 <= LB2D_shift_1;
       LB2D_shift_2 <= LB2D_shift_2;
       LB2D_shift_3 <= LB2D_shift_3;
       LB2D_shift_4 <= LB2D_shift_4;
       LB2D_shift_5 <= LB2D_shift_5;
       LB2D_shift_6 <= LB2D_shift_6;
       LB2D_shift_7 <= LB2D_shift_7;
       LB2D_shift_x <= LB2D_shift_x;
       LB2D_shift_y <= LB2D_shift_y;
       arg_0_TDATA <= arg_0_TDATA;
       arg_0_TVALID <= arg_0_TVALID;
       arg_1_TREADY <= arg_1_TREADY;
       gb_exit_it_1 <= gb_exit_it_1;
       gb_exit_it_2 <= gb_exit_it_2;
       gb_exit_it_3 <= gb_exit_it_3;
       gb_exit_it_4 <= gb_exit_it_4;
       gb_exit_it_5 <= gb_exit_it_5;
       gb_exit_it_6 <= gb_exit_it_6;
       gb_exit_it_7 <= gb_exit_it_7;
       gb_exit_it_8 <= gb_exit_it_8;
       gb_p_cnt <= gb_p_cnt;
       gb_pp_it_1 <= gb_pp_it_1;
       gb_pp_it_2 <= gb_pp_it_2;
       gb_pp_it_3 <= gb_pp_it_3;
       gb_pp_it_4 <= gb_pp_it_4;
       gb_pp_it_5 <= gb_pp_it_5;
       gb_pp_it_6 <= gb_pp_it_6;
       gb_pp_it_7 <= gb_pp_it_7;
       gb_pp_it_8 <= gb_pp_it_8;
       gb_pp_it_9 <= gb_pp_it_9;
       in_stream_buff_0 <= in_stream_buff_0;
       in_stream_buff_1 <= in_stream_buff_1;
       in_stream_empty <= in_stream_empty;
       in_stream_full <= in_stream_full;
       slice_stream_buff_0 <= slice_stream_buff_0;
       slice_stream_buff_1 <= slice_stream_buff_1;
       slice_stream_empty <= slice_stream_empty;
       slice_stream_full <= slice_stream_full;
       stencil_stream_buff_0 <= stencil_stream_buff_0;
       stencil_stream_buff_1 <= stencil_stream_buff_1;
       stencil_stream_empty <= stencil_stream_empty;
       stencil_stream_full <= stencil_stream_full;
   end
   else if(step) begin
       LB1D_buff <= n40;
       LB1D_in <= n46;
       LB1D_it_1 <= n50;
       LB1D_p_cnt <= n58;
       LB1D_uIn <= n63;
       LB2D_proc_w <= n73;
       LB2D_proc_x <= n80;
       LB2D_proc_y <= n89;
       LB2D_shift_0 <= n94;
       LB2D_shift_1 <= n99;
       LB2D_shift_2 <= n104;
       LB2D_shift_3 <= n109;
       LB2D_shift_4 <= n114;
       LB2D_shift_5 <= n119;
       LB2D_shift_6 <= n124;
       LB2D_shift_7 <= n131;
       LB2D_shift_x <= n137;
       LB2D_shift_y <= n147;
       arg_0_TDATA <= n155;
       arg_0_TVALID <= n162;
       arg_1_TREADY <= n171;
       gb_exit_it_1 <= n179;
       gb_exit_it_2 <= n184;
       gb_exit_it_3 <= n189;
       gb_exit_it_4 <= n194;
       gb_exit_it_5 <= n199;
       gb_exit_it_6 <= n204;
       gb_exit_it_7 <= n209;
       gb_exit_it_8 <= n214;
       gb_p_cnt <= n221;
       gb_pp_it_1 <= n226;
       gb_pp_it_2 <= n231;
       gb_pp_it_3 <= n236;
       gb_pp_it_4 <= n241;
       gb_pp_it_5 <= n246;
       gb_pp_it_6 <= n251;
       gb_pp_it_7 <= n256;
       gb_pp_it_8 <= n261;
       gb_pp_it_9 <= n266;
       in_stream_buff_0 <= n271;
       in_stream_buff_1 <= n276;
       in_stream_empty <= n283;
       in_stream_full <= n290;
       slice_stream_buff_0 <= n377;
       slice_stream_buff_1 <= n383;
       slice_stream_empty <= n390;
       slice_stream_full <= n398;
       stencil_stream_buff_0 <= n568;
       stencil_stream_buff_1 <= n573;
       stencil_stream_empty <= n581;
       stencil_stream_full <= n590;
       LB2D_proc_0 [ LB2D_proc_0_addr0 ] <= LB2D_proc_0_data0;
       LB2D_proc_1 [ LB2D_proc_1_addr0 ] <= LB2D_proc_1_data0;
       LB2D_proc_2 [ LB2D_proc_2_addr0 ] <= LB2D_proc_2_data0;
       LB2D_proc_3 [ LB2D_proc_3_addr0 ] <= LB2D_proc_3_data0;
       LB2D_proc_4 [ LB2D_proc_4_addr0 ] <= LB2D_proc_4_data0;
       LB2D_proc_5 [ LB2D_proc_5_addr0 ] <= LB2D_proc_5_data0;
       LB2D_proc_6 [ LB2D_proc_6_addr0 ] <= LB2D_proc_6_data0;
       LB2D_proc_7 [ LB2D_proc_7_addr0 ] <= LB2D_proc_7_data0;
   end
end
endmodule
