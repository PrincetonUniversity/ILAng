module GB(
arg_0_TREADY,
arg_1_TDATA,
arg_1_TVALID,
LB1D_buff,
LB2D_proc_w,
LB2D_proc_x,
LB2D_proc_y,
LB2D_shift_0,
LB2D_shift_1,
LB2D_shift_2,
LB2D_shift_3,
LB2D_shift_4,
LB2D_shift_5,
LB2D_shift_6,
LB2D_shift_7,
LB2D_shift_x,
LB2D_shift_y,
arg_0_TDATA,
arg_0_TVALID,
arg_1_TREADY,
in_stream_buff_0,
in_stream_buff_1,
in_stream_empty,
in_stream_full,
slice_stream_buff_0,
slice_stream_buff_1,
slice_stream_empty,
slice_stream_full,
stencil_stream_buff_0,
stencil_stream_buff_1,
stencil_stream_empty,
stencil_stream_full,
clk,rst,
step
);
input            arg_0_TREADY;
input      [7:0] arg_1_TDATA;
input            arg_1_TVALID;
input clk;
input rst;
input step;
output      [7:0] LB1D_buff;
output     [63:0] LB2D_proc_w;
output      [8:0] LB2D_proc_x;
output      [9:0] LB2D_proc_y;
output     [71:0] LB2D_shift_0;
output     [71:0] LB2D_shift_1;
output     [71:0] LB2D_shift_2;
output     [71:0] LB2D_shift_3;
output     [71:0] LB2D_shift_4;
output     [71:0] LB2D_shift_5;
output     [71:0] LB2D_shift_6;
output     [71:0] LB2D_shift_7;
output      [8:0] LB2D_shift_x;
output      [9:0] LB2D_shift_y;
output      [7:0] arg_0_TDATA;
output            arg_0_TVALID;
output            arg_1_TREADY;
output      [7:0] in_stream_buff_0;
output      [7:0] in_stream_buff_1;
output            in_stream_empty;
output            in_stream_full;
output     [71:0] slice_stream_buff_0;
output     [71:0] slice_stream_buff_1;
output            slice_stream_empty;
output            slice_stream_full;
output    [647:0] stencil_stream_buff_0;
output    [647:0] stencil_stream_buff_1;
output            stencil_stream_empty;
output            stencil_stream_full;
reg      [7:0] LB1D_buff;
reg     [63:0] LB2D_proc_w;
reg      [8:0] LB2D_proc_x;
reg      [9:0] LB2D_proc_y;
reg     [71:0] LB2D_shift_0;
reg     [71:0] LB2D_shift_1;
reg     [71:0] LB2D_shift_2;
reg     [71:0] LB2D_shift_3;
reg     [71:0] LB2D_shift_4;
reg     [71:0] LB2D_shift_5;
reg     [71:0] LB2D_shift_6;
reg     [71:0] LB2D_shift_7;
reg      [8:0] LB2D_shift_x;
reg      [9:0] LB2D_shift_y;
reg      [7:0] arg_0_TDATA;
reg            arg_0_TVALID;
reg            arg_1_TREADY;
reg      [7:0] in_stream_buff_0;
reg      [7:0] in_stream_buff_1;
reg            in_stream_empty;
reg            in_stream_full;
reg     [71:0] slice_stream_buff_0;
reg     [71:0] slice_stream_buff_1;
reg            slice_stream_empty;
reg            slice_stream_full;
reg    [647:0] stencil_stream_buff_0;
reg    [647:0] stencil_stream_buff_1;
reg            stencil_stream_empty;
reg            stencil_stream_full;
wire            arg_0_TREADY;
wire      [7:0] arg_1_TDATA;
wire            arg_1_TVALID;
wire            n0;
wire            n1;
wire            n2;
wire            n3;
wire            n4;
wire            n5;
wire            n6;
wire            n7;
wire            n8;
wire            n9;
wire            n10;
wire            n11;
wire            n12;
wire            n13;
wire            n14;
wire            n15;
wire            n16;
wire            n17;
wire            n18;
wire            n19;
wire            n20;
wire            n21;
wire            n22;
wire            n23;
wire            n24;
wire            n25;
wire      [7:0] n26;
wire      [7:0] n27;
wire      [7:0] n28;
wire      [7:0] n29;
wire      [7:0] n30;
wire      [7:0] n31;
wire            n32;
wire            n33;
wire     [63:0] n34;
wire     [63:0] n35;
wire     [63:0] n36;
wire     [63:0] n37;
wire     [63:0] n38;
wire     [63:0] n39;
wire     [63:0] n40;
wire     [63:0] n41;
wire     [63:0] n42;
wire      [8:0] n43;
wire      [8:0] n44;
wire      [8:0] n45;
wire      [8:0] n46;
wire      [8:0] n47;
wire      [8:0] n48;
wire      [8:0] n49;
wire      [8:0] n50;
wire            n51;
wire      [9:0] n52;
wire      [9:0] n53;
wire      [9:0] n54;
wire      [9:0] n55;
wire      [9:0] n56;
wire      [9:0] n57;
wire      [9:0] n58;
wire      [9:0] n59;
wire      [9:0] n60;
wire            n61;
wire     [71:0] n62;
wire     [71:0] n63;
wire     [71:0] n64;
wire     [71:0] n65;
wire     [71:0] n66;
wire     [71:0] n67;
wire     [71:0] n68;
wire     [71:0] n69;
wire     [71:0] n70;
wire     [71:0] n71;
wire     [71:0] n72;
wire     [71:0] n73;
wire     [71:0] n74;
wire     [71:0] n75;
wire     [71:0] n76;
wire     [71:0] n77;
wire     [71:0] n78;
wire     [71:0] n79;
wire     [71:0] n80;
wire     [71:0] n81;
wire     [71:0] n82;
wire     [71:0] n83;
wire     [71:0] n84;
wire     [71:0] n85;
wire     [71:0] n86;
wire     [71:0] n87;
wire     [71:0] n88;
wire     [71:0] n89;
wire     [71:0] n90;
wire     [71:0] n91;
wire     [71:0] n92;
wire     [71:0] n93;
wire     [71:0] n94;
wire     [71:0] n95;
wire     [71:0] n96;
wire     [71:0] n97;
wire     [71:0] n98;
wire     [71:0] n99;
wire     [71:0] n100;
wire     [71:0] n101;
wire     [71:0] n102;
wire     [71:0] n103;
wire     [71:0] n104;
wire     [71:0] n105;
wire     [71:0] n106;
wire     [71:0] n107;
wire     [71:0] n108;
wire     [71:0] n109;
wire     [71:0] n110;
wire            n111;
wire      [8:0] n112;
wire      [8:0] n113;
wire      [8:0] n114;
wire      [8:0] n115;
wire      [8:0] n116;
wire      [8:0] n117;
wire      [8:0] n118;
wire      [8:0] n119;
wire      [9:0] n120;
wire      [9:0] n121;
wire      [9:0] n122;
wire      [9:0] n123;
wire      [9:0] n124;
wire      [9:0] n125;
wire            n126;
wire    [647:0] n127;
wire      [7:0] n128;
wire      [7:0] n129;
wire      [7:0] n130;
wire      [7:0] n131;
wire      [7:0] n132;
wire      [7:0] n133;
wire      [7:0] n134;
wire            n135;
wire            n136;
wire            n137;
wire            n138;
wire            n139;
wire            n140;
wire            n141;
wire            n142;
wire            n143;
wire            n144;
wire            n145;
wire            n146;
wire      [7:0] n147;
wire      [7:0] n148;
wire      [7:0] n149;
wire      [7:0] n150;
wire      [7:0] n151;
wire      [7:0] n152;
wire      [7:0] n153;
wire      [7:0] n154;
wire      [7:0] n155;
wire      [7:0] n156;
wire      [7:0] n157;
wire      [7:0] n158;
wire            n159;
wire            n160;
wire            n161;
wire            n162;
wire            n163;
wire            n164;
wire            n165;
wire            n166;
wire            n167;
wire            n168;
wire            n169;
wire            n170;
wire            n171;
wire            n172;
wire            n173;
wire            n174;
wire      [7:0] n175;
wire            n176;
wire      [7:0] n177;
wire            n178;
wire      [7:0] n179;
wire            n180;
wire      [7:0] n181;
wire            n182;
wire      [7:0] n183;
wire            n184;
wire      [7:0] n185;
wire            n186;
wire      [7:0] n187;
wire            n188;
wire      [7:0] n189;
wire      [7:0] n190;
wire      [7:0] n191;
wire      [7:0] n192;
wire      [7:0] n193;
wire      [7:0] n194;
wire      [7:0] n195;
wire      [7:0] n196;
wire      [7:0] n197;
wire      [7:0] n198;
wire      [7:0] n199;
wire      [7:0] n200;
wire      [7:0] n201;
wire      [7:0] n202;
wire      [7:0] n203;
wire      [7:0] n204;
wire      [7:0] n205;
wire      [7:0] n206;
wire      [7:0] n207;
wire      [7:0] n208;
wire      [7:0] n209;
wire      [7:0] n210;
wire      [7:0] n211;
wire      [7:0] n212;
wire      [7:0] n213;
wire      [7:0] n214;
wire      [7:0] n215;
wire      [7:0] n216;
wire      [7:0] n217;
wire      [7:0] n218;
wire      [7:0] n219;
wire      [7:0] n220;
wire      [7:0] n221;
wire      [7:0] n222;
wire      [7:0] n223;
wire      [7:0] n224;
wire      [7:0] n225;
wire      [7:0] n226;
wire      [7:0] n227;
wire      [7:0] n228;
wire      [7:0] n229;
wire      [7:0] n230;
wire      [7:0] n231;
wire      [7:0] n232;
wire      [7:0] n233;
wire      [7:0] n234;
wire      [7:0] n235;
wire      [7:0] n236;
wire      [7:0] n237;
wire      [7:0] n238;
wire      [7:0] n239;
wire      [7:0] n240;
wire      [7:0] n241;
wire      [7:0] n242;
wire      [7:0] n243;
wire      [7:0] n244;
wire      [7:0] n245;
wire      [7:0] n246;
wire     [15:0] n247;
wire     [23:0] n248;
wire     [31:0] n249;
wire     [39:0] n250;
wire     [47:0] n251;
wire     [55:0] n252;
wire     [63:0] n253;
wire     [71:0] n254;
wire     [71:0] n255;
wire     [71:0] n256;
wire     [71:0] n257;
wire     [71:0] n258;
wire     [71:0] n259;
wire     [71:0] n260;
wire     [71:0] n261;
wire     [71:0] n262;
wire     [71:0] n263;
wire     [71:0] n264;
wire     [71:0] n265;
wire     [71:0] n266;
wire     [71:0] n267;
wire     [71:0] n268;
wire            n269;
wire            n270;
wire            n271;
wire            n272;
wire            n273;
wire            n274;
wire            n275;
wire            n276;
wire            n277;
wire            n278;
wire            n279;
wire            n280;
wire            n281;
wire            n282;
wire            n283;
wire            n284;
wire            n285;
wire            n286;
wire      [7:0] n287;
wire      [7:0] n288;
wire      [7:0] n289;
wire      [7:0] n290;
wire      [7:0] n291;
wire      [7:0] n292;
wire      [7:0] n293;
wire      [7:0] n294;
wire      [7:0] n295;
wire     [15:0] n296;
wire     [23:0] n297;
wire     [31:0] n298;
wire     [39:0] n299;
wire     [47:0] n300;
wire     [55:0] n301;
wire     [63:0] n302;
wire     [71:0] n303;
wire      [7:0] n304;
wire      [7:0] n305;
wire      [7:0] n306;
wire      [7:0] n307;
wire      [7:0] n308;
wire      [7:0] n309;
wire      [7:0] n310;
wire      [7:0] n311;
wire      [7:0] n312;
wire     [15:0] n313;
wire     [23:0] n314;
wire     [31:0] n315;
wire     [39:0] n316;
wire     [47:0] n317;
wire     [55:0] n318;
wire     [63:0] n319;
wire     [71:0] n320;
wire      [7:0] n321;
wire      [7:0] n322;
wire      [7:0] n323;
wire      [7:0] n324;
wire      [7:0] n325;
wire      [7:0] n326;
wire      [7:0] n327;
wire      [7:0] n328;
wire      [7:0] n329;
wire     [15:0] n330;
wire     [23:0] n331;
wire     [31:0] n332;
wire     [39:0] n333;
wire     [47:0] n334;
wire     [55:0] n335;
wire     [63:0] n336;
wire     [71:0] n337;
wire      [7:0] n338;
wire      [7:0] n339;
wire      [7:0] n340;
wire      [7:0] n341;
wire      [7:0] n342;
wire      [7:0] n343;
wire      [7:0] n344;
wire      [7:0] n345;
wire      [7:0] n346;
wire     [15:0] n347;
wire     [23:0] n348;
wire     [31:0] n349;
wire     [39:0] n350;
wire     [47:0] n351;
wire     [55:0] n352;
wire     [63:0] n353;
wire     [71:0] n354;
wire      [7:0] n355;
wire      [7:0] n356;
wire      [7:0] n357;
wire      [7:0] n358;
wire      [7:0] n359;
wire      [7:0] n360;
wire      [7:0] n361;
wire      [7:0] n362;
wire      [7:0] n363;
wire     [15:0] n364;
wire     [23:0] n365;
wire     [31:0] n366;
wire     [39:0] n367;
wire     [47:0] n368;
wire     [55:0] n369;
wire     [63:0] n370;
wire     [71:0] n371;
wire      [7:0] n372;
wire      [7:0] n373;
wire      [7:0] n374;
wire      [7:0] n375;
wire      [7:0] n376;
wire      [7:0] n377;
wire      [7:0] n378;
wire      [7:0] n379;
wire      [7:0] n380;
wire     [15:0] n381;
wire     [23:0] n382;
wire     [31:0] n383;
wire     [39:0] n384;
wire     [47:0] n385;
wire     [55:0] n386;
wire     [63:0] n387;
wire     [71:0] n388;
wire      [7:0] n389;
wire      [7:0] n390;
wire      [7:0] n391;
wire      [7:0] n392;
wire      [7:0] n393;
wire      [7:0] n394;
wire      [7:0] n395;
wire      [7:0] n396;
wire      [7:0] n397;
wire     [15:0] n398;
wire     [23:0] n399;
wire     [31:0] n400;
wire     [39:0] n401;
wire     [47:0] n402;
wire     [55:0] n403;
wire     [63:0] n404;
wire     [71:0] n405;
wire      [7:0] n406;
wire      [7:0] n407;
wire      [7:0] n408;
wire      [7:0] n409;
wire      [7:0] n410;
wire      [7:0] n411;
wire      [7:0] n412;
wire      [7:0] n413;
wire      [7:0] n414;
wire     [15:0] n415;
wire     [23:0] n416;
wire     [31:0] n417;
wire     [39:0] n418;
wire     [47:0] n419;
wire     [55:0] n420;
wire     [63:0] n421;
wire     [71:0] n422;
wire      [7:0] n423;
wire      [7:0] n424;
wire      [7:0] n425;
wire      [7:0] n426;
wire      [7:0] n427;
wire      [7:0] n428;
wire      [7:0] n429;
wire      [7:0] n430;
wire      [7:0] n431;
wire     [15:0] n432;
wire     [23:0] n433;
wire     [31:0] n434;
wire     [39:0] n435;
wire     [47:0] n436;
wire     [55:0] n437;
wire     [63:0] n438;
wire     [71:0] n439;
wire    [143:0] n440;
wire    [215:0] n441;
wire    [287:0] n442;
wire    [359:0] n443;
wire    [431:0] n444;
wire    [503:0] n445;
wire    [575:0] n446;
wire    [647:0] n447;
wire    [647:0] n448;
wire    [647:0] n449;
wire    [647:0] n450;
wire    [647:0] n451;
wire    [647:0] n452;
wire    [647:0] n453;
wire    [647:0] n454;
wire    [647:0] n455;
wire    [647:0] n456;
wire    [647:0] n457;
wire    [647:0] n458;
wire    [647:0] n459;
wire    [647:0] n460;
wire            n461;
wire            n462;
wire            n463;
wire            n464;
wire            n465;
wire            n466;
wire            n467;
wire            n468;
wire            n469;
wire            n470;
wire            n471;
wire            n472;
wire            n473;
wire            n474;
wire            n475;
wire            n476;
wire            n477;
wire      [8:0] LB2D_proc_0_addr0;
wire      [7:0] LB2D_proc_0_data0;
wire            n478;
wire            n479;
wire            n480;
wire            n481;
wire            n482;
wire            n483;
wire            n484;
wire            n485;
wire            n486;
wire            n487;
wire            n488;
wire            n489;
wire            n490;
wire            n491;
wire            n492;
wire            n493;
wire            n494;
wire            n495;
wire            n496;
wire      [8:0] LB2D_proc_1_addr0;
wire      [7:0] LB2D_proc_1_data0;
wire            n497;
wire            n498;
wire            n499;
wire      [8:0] LB2D_proc_2_addr0;
wire      [7:0] LB2D_proc_2_data0;
wire            n500;
wire            n501;
wire            n502;
wire      [8:0] LB2D_proc_3_addr0;
wire      [7:0] LB2D_proc_3_data0;
wire            n503;
wire            n504;
wire            n505;
wire      [8:0] LB2D_proc_4_addr0;
wire      [7:0] LB2D_proc_4_data0;
wire            n506;
wire            n507;
wire            n508;
wire      [8:0] LB2D_proc_5_addr0;
wire      [7:0] LB2D_proc_5_data0;
wire            n509;
wire            n510;
wire            n511;
wire      [8:0] LB2D_proc_6_addr0;
wire      [7:0] LB2D_proc_6_data0;
wire            n512;
wire            n513;
wire            n514;
wire      [8:0] LB2D_proc_7_addr0;
wire      [7:0] LB2D_proc_7_data0;
wire            n515;
wire            n516;
wire            n517;
wire            n518;
reg      [7:0] LB2D_proc_0[511:0];
reg      [7:0] LB2D_proc_1[511:0];
reg      [7:0] LB2D_proc_2[511:0];
reg      [7:0] LB2D_proc_3[511:0];
reg      [7:0] LB2D_proc_4[511:0];
reg      [7:0] LB2D_proc_5[511:0];
reg      [7:0] LB2D_proc_6[511:0];
reg      [7:0] LB2D_proc_7[511:0];
wire clk;
wire rst;
wire step;
assign n0 =  ( arg_0_TREADY ) == ( 1'd1 )  ;
assign n1 =  ( arg_0_TVALID ) == ( 1'd1 )  ;
assign n2 =  ( n0 ) & ( n1 )  ;
assign n3 =  ( arg_1_TVALID ) == ( 1'd0 )  ;
assign n4 =  ( n2 ) & ( n3 )  ;
assign n5 =  ( arg_1_TREADY ) == ( 1'd1 )  ;
assign n6 =  ( arg_1_TVALID ) == ( 1'd1 )  ;
assign n7 =  ( n5 ) & ( n6 )  ;
assign n8 =  ( arg_0_TREADY ) == ( 1'd0 )  ;
assign n9 =  ( n7 ) & ( n8 )  ;
assign n10 =  ( stencil_stream_empty ) == ( 1'd0 )  ;
assign n11 =  ( arg_0_TVALID ) == ( 1'd0 )  ;
assign n12 =  ( n10 ) & ( n11 )  ;
assign n13 =  ( slice_stream_empty ) == ( 1'd0 )  ;
assign n14 =  ( stencil_stream_full ) == ( 1'd0 )  ;
assign n15 =  ( LB2D_shift_x ) < ( 9'd8 )  ;
assign n16 =  ( n14 ) | ( n15 )  ;
assign n17 =  ( n13 ) & ( n16 )  ;
assign n18 =  ( in_stream_empty ) == ( 1'd0 )  ;
assign n19 =  ( slice_stream_full ) == ( 1'd0 )  ;
assign n20 =  ( LB2D_proc_y ) < ( 10'd8 )  ;
assign n21 =  ( n19 ) | ( n20 )  ;
assign n22 =  ( n18 ) & ( n21 )  ;
assign n23 =  ( arg_1_TREADY ) == ( 1'd0 )  ;
assign n24 =  ( in_stream_full ) == ( 1'd0 )  ;
assign n25 =  ( n23 ) & ( n24 )  ;
assign n26 =  ( n25 ) ? ( LB1D_buff ) : ( LB1D_buff ) ;
assign n27 =  ( n22 ) ? ( LB1D_buff ) : ( n26 ) ;
assign n28 =  ( n17 ) ? ( LB1D_buff ) : ( n27 ) ;
assign n29 =  ( n12 ) ? ( LB1D_buff ) : ( n28 ) ;
assign n30 =  ( n9 ) ? ( arg_1_TDATA ) : ( n29 ) ;
assign n31 =  ( n4 ) ? ( arg_1_TDATA ) : ( n30 ) ;
assign n32 =  ( LB2D_proc_w ) < ( 64'd7 )  ;
assign n33 =  ( LB2D_proc_x ) < ( 9'd487 )  ;
assign n34 =  ( LB2D_proc_w ) + ( 64'd1 )  ;
assign n35 =  ( n33 ) ? ( LB2D_proc_w ) : ( n34 ) ;
assign n36 =  ( n32 ) ? ( n35 ) : ( 64'd0 ) ;
assign n37 =  ( n25 ) ? ( LB2D_proc_w ) : ( LB2D_proc_w ) ;
assign n38 =  ( n22 ) ? ( n36 ) : ( n37 ) ;
assign n39 =  ( n17 ) ? ( LB2D_proc_w ) : ( n38 ) ;
assign n40 =  ( n12 ) ? ( LB2D_proc_w ) : ( n39 ) ;
assign n41 =  ( n9 ) ? ( LB2D_proc_w ) : ( n40 ) ;
assign n42 =  ( n4 ) ? ( LB2D_proc_w ) : ( n41 ) ;
assign n43 =  ( LB2D_proc_x ) + ( 9'd1 )  ;
assign n44 =  ( n33 ) ? ( n43 ) : ( 9'd0 ) ;
assign n45 =  ( n25 ) ? ( LB2D_proc_x ) : ( LB2D_proc_x ) ;
assign n46 =  ( n22 ) ? ( n44 ) : ( n45 ) ;
assign n47 =  ( n17 ) ? ( LB2D_proc_x ) : ( n46 ) ;
assign n48 =  ( n12 ) ? ( LB2D_proc_x ) : ( n47 ) ;
assign n49 =  ( n9 ) ? ( LB2D_proc_x ) : ( n48 ) ;
assign n50 =  ( n4 ) ? ( LB2D_proc_x ) : ( n49 ) ;
assign n51 =  ( LB2D_proc_y ) < ( 10'd487 )  ;
assign n52 =  ( LB2D_proc_y ) + ( 10'd1 )  ;
assign n53 =  ( n33 ) ? ( LB2D_proc_y ) : ( n52 ) ;
assign n54 =  ( n51 ) ? ( n53 ) : ( 10'd487 ) ;
assign n55 =  ( n25 ) ? ( LB2D_proc_y ) : ( LB2D_proc_y ) ;
assign n56 =  ( n22 ) ? ( n54 ) : ( n55 ) ;
assign n57 =  ( n17 ) ? ( LB2D_proc_y ) : ( n56 ) ;
assign n58 =  ( n12 ) ? ( LB2D_proc_y ) : ( n57 ) ;
assign n59 =  ( n9 ) ? ( LB2D_proc_y ) : ( n58 ) ;
assign n60 =  ( n4 ) ? ( LB2D_proc_y ) : ( n59 ) ;
assign n61 =  ( slice_stream_full ) == ( 1'd1 )  ;
assign n62 =  ( n61 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n63 =  ( n25 ) ? ( LB2D_shift_0 ) : ( LB2D_shift_0 ) ;
assign n64 =  ( n22 ) ? ( LB2D_shift_0 ) : ( n63 ) ;
assign n65 =  ( n17 ) ? ( n62 ) : ( n64 ) ;
assign n66 =  ( n12 ) ? ( LB2D_shift_0 ) : ( n65 ) ;
assign n67 =  ( n9 ) ? ( LB2D_shift_0 ) : ( n66 ) ;
assign n68 =  ( n4 ) ? ( LB2D_shift_0 ) : ( n67 ) ;
assign n69 =  ( n25 ) ? ( LB2D_shift_1 ) : ( LB2D_shift_1 ) ;
assign n70 =  ( n22 ) ? ( LB2D_shift_1 ) : ( n69 ) ;
assign n71 =  ( n17 ) ? ( LB2D_shift_0 ) : ( n70 ) ;
assign n72 =  ( n12 ) ? ( LB2D_shift_1 ) : ( n71 ) ;
assign n73 =  ( n9 ) ? ( LB2D_shift_1 ) : ( n72 ) ;
assign n74 =  ( n4 ) ? ( LB2D_shift_1 ) : ( n73 ) ;
assign n75 =  ( n25 ) ? ( LB2D_shift_2 ) : ( LB2D_shift_2 ) ;
assign n76 =  ( n22 ) ? ( LB2D_shift_2 ) : ( n75 ) ;
assign n77 =  ( n17 ) ? ( LB2D_shift_1 ) : ( n76 ) ;
assign n78 =  ( n12 ) ? ( LB2D_shift_2 ) : ( n77 ) ;
assign n79 =  ( n9 ) ? ( LB2D_shift_2 ) : ( n78 ) ;
assign n80 =  ( n4 ) ? ( LB2D_shift_2 ) : ( n79 ) ;
assign n81 =  ( n25 ) ? ( LB2D_shift_3 ) : ( LB2D_shift_3 ) ;
assign n82 =  ( n22 ) ? ( LB2D_shift_3 ) : ( n81 ) ;
assign n83 =  ( n17 ) ? ( LB2D_shift_2 ) : ( n82 ) ;
assign n84 =  ( n12 ) ? ( LB2D_shift_3 ) : ( n83 ) ;
assign n85 =  ( n9 ) ? ( LB2D_shift_3 ) : ( n84 ) ;
assign n86 =  ( n4 ) ? ( LB2D_shift_3 ) : ( n85 ) ;
assign n87 =  ( n25 ) ? ( LB2D_shift_4 ) : ( LB2D_shift_4 ) ;
assign n88 =  ( n22 ) ? ( LB2D_shift_4 ) : ( n87 ) ;
assign n89 =  ( n17 ) ? ( LB2D_shift_3 ) : ( n88 ) ;
assign n90 =  ( n12 ) ? ( LB2D_shift_4 ) : ( n89 ) ;
assign n91 =  ( n9 ) ? ( LB2D_shift_4 ) : ( n90 ) ;
assign n92 =  ( n4 ) ? ( LB2D_shift_4 ) : ( n91 ) ;
assign n93 =  ( n25 ) ? ( LB2D_shift_5 ) : ( LB2D_shift_5 ) ;
assign n94 =  ( n22 ) ? ( LB2D_shift_5 ) : ( n93 ) ;
assign n95 =  ( n17 ) ? ( LB2D_shift_4 ) : ( n94 ) ;
assign n96 =  ( n12 ) ? ( LB2D_shift_5 ) : ( n95 ) ;
assign n97 =  ( n9 ) ? ( LB2D_shift_5 ) : ( n96 ) ;
assign n98 =  ( n4 ) ? ( LB2D_shift_5 ) : ( n97 ) ;
assign n99 =  ( n25 ) ? ( LB2D_shift_6 ) : ( LB2D_shift_6 ) ;
assign n100 =  ( n22 ) ? ( LB2D_shift_6 ) : ( n99 ) ;
assign n101 =  ( n17 ) ? ( LB2D_shift_5 ) : ( n100 ) ;
assign n102 =  ( n12 ) ? ( LB2D_shift_6 ) : ( n101 ) ;
assign n103 =  ( n9 ) ? ( LB2D_shift_6 ) : ( n102 ) ;
assign n104 =  ( n4 ) ? ( LB2D_shift_6 ) : ( n103 ) ;
assign n105 =  ( n25 ) ? ( LB2D_shift_7 ) : ( LB2D_shift_7 ) ;
assign n106 =  ( n22 ) ? ( LB2D_shift_7 ) : ( n105 ) ;
assign n107 =  ( n17 ) ? ( LB2D_shift_6 ) : ( n106 ) ;
assign n108 =  ( n12 ) ? ( LB2D_shift_7 ) : ( n107 ) ;
assign n109 =  ( n9 ) ? ( LB2D_shift_7 ) : ( n108 ) ;
assign n110 =  ( n4 ) ? ( LB2D_shift_7 ) : ( n109 ) ;
assign n111 =  ( LB2D_shift_x ) < ( 9'd487 )  ;
assign n112 =  ( LB2D_shift_x ) + ( 9'd1 )  ;
assign n113 =  ( n111 ) ? ( n112 ) : ( 9'd0 ) ;
assign n114 =  ( n25 ) ? ( LB2D_shift_x ) : ( LB2D_shift_x ) ;
assign n115 =  ( n22 ) ? ( LB2D_shift_x ) : ( n114 ) ;
assign n116 =  ( n17 ) ? ( n113 ) : ( n115 ) ;
assign n117 =  ( n12 ) ? ( LB2D_shift_x ) : ( n116 ) ;
assign n118 =  ( n9 ) ? ( LB2D_shift_x ) : ( n117 ) ;
assign n119 =  ( n4 ) ? ( LB2D_shift_x ) : ( n118 ) ;
assign n120 =  ( n25 ) ? ( LB2D_shift_y ) : ( LB2D_shift_y ) ;
assign n121 =  ( n22 ) ? ( LB2D_shift_y ) : ( n120 ) ;
assign n122 =  ( n17 ) ? ( LB2D_shift_y ) : ( n121 ) ;
assign n123 =  ( n12 ) ? ( LB2D_shift_y ) : ( n122 ) ;
assign n124 =  ( n9 ) ? ( LB2D_shift_y ) : ( n123 ) ;
assign n125 =  ( n4 ) ? ( LB2D_shift_y ) : ( n124 ) ;
assign n126 =  ( stencil_stream_full ) == ( 1'd1 )  ;
assign n127 =  ( n126 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_0 ) ;
//assign n128 = gb_fun(n127) ;
gb_fun gb_fun_U (
    .stencil (n127),
    .result (n128)
);


assign n129 =  ( n25 ) ? ( arg_0_TDATA ) : ( arg_0_TDATA ) ;
assign n130 =  ( n22 ) ? ( arg_0_TDATA ) : ( n129 ) ;
assign n131 =  ( n17 ) ? ( arg_0_TDATA ) : ( n130 ) ;
assign n132 =  ( n12 ) ? ( n128 ) : ( n131 ) ;
assign n133 =  ( n9 ) ? ( arg_0_TDATA ) : ( n132 ) ;
assign n134 =  ( n4 ) ? ( arg_0_TDATA ) : ( n133 ) ;
assign n135 =  ( n25 ) ? ( arg_0_TVALID ) : ( arg_0_TVALID ) ;
assign n136 =  ( n22 ) ? ( arg_0_TVALID ) : ( n135 ) ;
assign n137 =  ( n17 ) ? ( arg_0_TVALID ) : ( n136 ) ;
assign n138 =  ( n12 ) ? ( 1'd1 ) : ( n137 ) ;
assign n139 =  ( n9 ) ? ( arg_0_TVALID ) : ( n138 ) ;
assign n140 =  ( n4 ) ? ( 1'd0 ) : ( n139 ) ;
assign n141 =  ( n25 ) ? ( 1'd1 ) : ( arg_1_TREADY ) ;
assign n142 =  ( n22 ) ? ( arg_1_TREADY ) : ( n141 ) ;
assign n143 =  ( n17 ) ? ( arg_1_TREADY ) : ( n142 ) ;
assign n144 =  ( n12 ) ? ( arg_1_TREADY ) : ( n143 ) ;
assign n145 =  ( n9 ) ? ( 1'd0 ) : ( n144 ) ;
assign n146 =  ( n4 ) ? ( 1'd0 ) : ( n145 ) ;
assign n147 =  ( n25 ) ? ( LB1D_buff ) : ( in_stream_buff_0 ) ;
assign n148 =  ( n22 ) ? ( in_stream_buff_0 ) : ( n147 ) ;
assign n149 =  ( n17 ) ? ( in_stream_buff_0 ) : ( n148 ) ;
assign n150 =  ( n12 ) ? ( in_stream_buff_0 ) : ( n149 ) ;
assign n151 =  ( n9 ) ? ( in_stream_buff_0 ) : ( n150 ) ;
assign n152 =  ( n4 ) ? ( in_stream_buff_0 ) : ( n151 ) ;
assign n153 =  ( n25 ) ? ( in_stream_buff_0 ) : ( in_stream_buff_1 ) ;
assign n154 =  ( n22 ) ? ( in_stream_buff_1 ) : ( n153 ) ;
assign n155 =  ( n17 ) ? ( in_stream_buff_1 ) : ( n154 ) ;
assign n156 =  ( n12 ) ? ( in_stream_buff_1 ) : ( n155 ) ;
assign n157 =  ( n9 ) ? ( in_stream_buff_1 ) : ( n156 ) ;
assign n158 =  ( n4 ) ? ( in_stream_buff_1 ) : ( n157 ) ;
assign n159 =  ( in_stream_full ) == ( 1'd1 )  ;
assign n160 =  ( n159 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n161 =  ( n25 ) ? ( 1'd0 ) : ( in_stream_empty ) ;
assign n162 =  ( n22 ) ? ( n160 ) : ( n161 ) ;
assign n163 =  ( n17 ) ? ( in_stream_empty ) : ( n162 ) ;
assign n164 =  ( n12 ) ? ( in_stream_empty ) : ( n163 ) ;
assign n165 =  ( n9 ) ? ( in_stream_empty ) : ( n164 ) ;
assign n166 =  ( n4 ) ? ( in_stream_empty ) : ( n165 ) ;
assign n167 =  ( in_stream_empty ) == ( 1'd1 )  ;
assign n168 =  ( n167 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n169 =  ( n25 ) ? ( n168 ) : ( in_stream_full ) ;
assign n170 =  ( n22 ) ? ( 1'd0 ) : ( n169 ) ;
assign n171 =  ( n17 ) ? ( in_stream_full ) : ( n170 ) ;
assign n172 =  ( n12 ) ? ( in_stream_full ) : ( n171 ) ;
assign n173 =  ( n9 ) ? ( in_stream_full ) : ( n172 ) ;
assign n174 =  ( n4 ) ? ( in_stream_full ) : ( n173 ) ;
assign n175 =  ( n159 ) ? ( in_stream_buff_1 ) : ( in_stream_buff_0 ) ;
assign n176 =  ( LB2D_proc_w ) == ( 64'd0 )  ;
assign n177 =  (  LB2D_proc_7 [ LB2D_proc_x ] )  ;
assign n178 =  ( LB2D_proc_w ) == ( 64'd1 )  ;
assign n179 =  (  LB2D_proc_0 [ LB2D_proc_x ] )  ;
assign n180 =  ( LB2D_proc_w ) == ( 64'd2 )  ;
assign n181 =  (  LB2D_proc_1 [ LB2D_proc_x ] )  ;
assign n182 =  ( LB2D_proc_w ) == ( 64'd3 )  ;
assign n183 =  (  LB2D_proc_2 [ LB2D_proc_x ] )  ;
assign n184 =  ( LB2D_proc_w ) == ( 64'd4 )  ;
assign n185 =  (  LB2D_proc_3 [ LB2D_proc_x ] )  ;
assign n186 =  ( LB2D_proc_w ) == ( 64'd5 )  ;
assign n187 =  (  LB2D_proc_4 [ LB2D_proc_x ] )  ;
assign n188 =  ( LB2D_proc_w ) == ( 64'd6 )  ;
assign n189 =  (  LB2D_proc_5 [ LB2D_proc_x ] )  ;
assign n190 =  (  LB2D_proc_6 [ LB2D_proc_x ] )  ;
assign n191 =  ( n188 ) ? ( n189 ) : ( n190 ) ;
assign n192 =  ( n186 ) ? ( n187 ) : ( n191 ) ;
assign n193 =  ( n184 ) ? ( n185 ) : ( n192 ) ;
assign n194 =  ( n182 ) ? ( n183 ) : ( n193 ) ;
assign n195 =  ( n180 ) ? ( n181 ) : ( n194 ) ;
assign n196 =  ( n178 ) ? ( n179 ) : ( n195 ) ;
assign n197 =  ( n176 ) ? ( n177 ) : ( n196 ) ;
assign n198 =  ( n188 ) ? ( n187 ) : ( n189 ) ;
assign n199 =  ( n186 ) ? ( n185 ) : ( n198 ) ;
assign n200 =  ( n184 ) ? ( n183 ) : ( n199 ) ;
assign n201 =  ( n182 ) ? ( n181 ) : ( n200 ) ;
assign n202 =  ( n180 ) ? ( n179 ) : ( n201 ) ;
assign n203 =  ( n178 ) ? ( n177 ) : ( n202 ) ;
assign n204 =  ( n176 ) ? ( n190 ) : ( n203 ) ;
assign n205 =  ( n188 ) ? ( n185 ) : ( n187 ) ;
assign n206 =  ( n186 ) ? ( n183 ) : ( n205 ) ;
assign n207 =  ( n184 ) ? ( n181 ) : ( n206 ) ;
assign n208 =  ( n182 ) ? ( n179 ) : ( n207 ) ;
assign n209 =  ( n180 ) ? ( n177 ) : ( n208 ) ;
assign n210 =  ( n178 ) ? ( n190 ) : ( n209 ) ;
assign n211 =  ( n176 ) ? ( n189 ) : ( n210 ) ;
assign n212 =  ( n188 ) ? ( n183 ) : ( n185 ) ;
assign n213 =  ( n186 ) ? ( n181 ) : ( n212 ) ;
assign n214 =  ( n184 ) ? ( n179 ) : ( n213 ) ;
assign n215 =  ( n182 ) ? ( n177 ) : ( n214 ) ;
assign n216 =  ( n180 ) ? ( n190 ) : ( n215 ) ;
assign n217 =  ( n178 ) ? ( n189 ) : ( n216 ) ;
assign n218 =  ( n176 ) ? ( n187 ) : ( n217 ) ;
assign n219 =  ( n188 ) ? ( n181 ) : ( n183 ) ;
assign n220 =  ( n186 ) ? ( n179 ) : ( n219 ) ;
assign n221 =  ( n184 ) ? ( n177 ) : ( n220 ) ;
assign n222 =  ( n182 ) ? ( n190 ) : ( n221 ) ;
assign n223 =  ( n180 ) ? ( n189 ) : ( n222 ) ;
assign n224 =  ( n178 ) ? ( n187 ) : ( n223 ) ;
assign n225 =  ( n176 ) ? ( n185 ) : ( n224 ) ;
assign n226 =  ( n188 ) ? ( n179 ) : ( n181 ) ;
assign n227 =  ( n186 ) ? ( n177 ) : ( n226 ) ;
assign n228 =  ( n184 ) ? ( n190 ) : ( n227 ) ;
assign n229 =  ( n182 ) ? ( n189 ) : ( n228 ) ;
assign n230 =  ( n180 ) ? ( n187 ) : ( n229 ) ;
assign n231 =  ( n178 ) ? ( n185 ) : ( n230 ) ;
assign n232 =  ( n176 ) ? ( n183 ) : ( n231 ) ;
assign n233 =  ( n188 ) ? ( n177 ) : ( n179 ) ;
assign n234 =  ( n186 ) ? ( n190 ) : ( n233 ) ;
assign n235 =  ( n184 ) ? ( n189 ) : ( n234 ) ;
assign n236 =  ( n182 ) ? ( n187 ) : ( n235 ) ;
assign n237 =  ( n180 ) ? ( n185 ) : ( n236 ) ;
assign n238 =  ( n178 ) ? ( n183 ) : ( n237 ) ;
assign n239 =  ( n176 ) ? ( n181 ) : ( n238 ) ;
assign n240 =  ( n188 ) ? ( n190 ) : ( n177 ) ;
assign n241 =  ( n186 ) ? ( n189 ) : ( n240 ) ;
assign n242 =  ( n184 ) ? ( n187 ) : ( n241 ) ;
assign n243 =  ( n182 ) ? ( n185 ) : ( n242 ) ;
assign n244 =  ( n180 ) ? ( n183 ) : ( n243 ) ;
assign n245 =  ( n178 ) ? ( n181 ) : ( n244 ) ;
assign n246 =  ( n176 ) ? ( n179 ) : ( n245 ) ;
assign n247 =  { ( n239 ) , ( n246 ) }  ;
assign n248 =  { ( n232 ) , ( n247 ) }  ;
assign n249 =  { ( n225 ) , ( n248 ) }  ;
assign n250 =  { ( n218 ) , ( n249 ) }  ;
assign n251 =  { ( n211 ) , ( n250 ) }  ;
assign n252 =  { ( n204 ) , ( n251 ) }  ;
assign n253 =  { ( n197 ) , ( n252 ) }  ;
assign n254 =  { ( n175 ) , ( n253 ) }  ;
assign n255 =  ( n20 ) ? ( slice_stream_buff_0 ) : ( n254 ) ;
assign n256 =  ( n25 ) ? ( slice_stream_buff_0 ) : ( slice_stream_buff_0 ) ;
assign n257 =  ( n22 ) ? ( n255 ) : ( n256 ) ;
assign n258 =  ( n17 ) ? ( slice_stream_buff_0 ) : ( n257 ) ;
assign n259 =  ( n12 ) ? ( slice_stream_buff_0 ) : ( n258 ) ;
assign n260 =  ( n9 ) ? ( slice_stream_buff_0 ) : ( n259 ) ;
assign n261 =  ( n4 ) ? ( slice_stream_buff_0 ) : ( n260 ) ;
assign n262 =  ( n20 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n263 =  ( n25 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_1 ) ;
assign n264 =  ( n22 ) ? ( n262 ) : ( n263 ) ;
assign n265 =  ( n17 ) ? ( slice_stream_buff_1 ) : ( n264 ) ;
assign n266 =  ( n12 ) ? ( slice_stream_buff_1 ) : ( n265 ) ;
assign n267 =  ( n9 ) ? ( slice_stream_buff_1 ) : ( n266 ) ;
assign n268 =  ( n4 ) ? ( slice_stream_buff_1 ) : ( n267 ) ;
assign n269 =  ( n61 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n270 =  ( n20 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n271 =  ( n25 ) ? ( slice_stream_empty ) : ( slice_stream_empty ) ;
assign n272 =  ( n22 ) ? ( n270 ) : ( n271 ) ;
assign n273 =  ( n17 ) ? ( n269 ) : ( n272 ) ;
assign n274 =  ( n12 ) ? ( slice_stream_empty ) : ( n273 ) ;
assign n275 =  ( n9 ) ? ( slice_stream_empty ) : ( n274 ) ;
assign n276 =  ( n4 ) ? ( slice_stream_empty ) : ( n275 ) ;
assign n277 =  ( slice_stream_empty ) == ( 1'd1 )  ;
assign n278 =  ( n277 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n279 =  ( n20 ) ? ( 1'd0 ) : ( n278 ) ;
assign n280 =  ( n25 ) ? ( slice_stream_full ) : ( slice_stream_full ) ;
assign n281 =  ( n22 ) ? ( n279 ) : ( n280 ) ;
assign n282 =  ( n17 ) ? ( 1'd0 ) : ( n281 ) ;
assign n283 =  ( n12 ) ? ( slice_stream_full ) : ( n282 ) ;
assign n284 =  ( n9 ) ? ( slice_stream_full ) : ( n283 ) ;
assign n285 =  ( n4 ) ? ( slice_stream_full ) : ( n284 ) ;
assign n286 =  ( LB2D_shift_x ) >= ( 9'd8 )  ;
assign n287 = n62[71:64] ;
assign n288 = LB2D_shift_0[71:64] ;
assign n289 = LB2D_shift_1[71:64] ;
assign n290 = LB2D_shift_2[71:64] ;
assign n291 = LB2D_shift_3[71:64] ;
assign n292 = LB2D_shift_4[71:64] ;
assign n293 = LB2D_shift_5[71:64] ;
assign n294 = LB2D_shift_6[71:64] ;
assign n295 = LB2D_shift_7[71:64] ;
assign n296 =  { ( n294 ) , ( n295 ) }  ;
assign n297 =  { ( n293 ) , ( n296 ) }  ;
assign n298 =  { ( n292 ) , ( n297 ) }  ;
assign n299 =  { ( n291 ) , ( n298 ) }  ;
assign n300 =  { ( n290 ) , ( n299 ) }  ;
assign n301 =  { ( n289 ) , ( n300 ) }  ;
assign n302 =  { ( n288 ) , ( n301 ) }  ;
assign n303 =  { ( n287 ) , ( n302 ) }  ;
assign n304 = n62[63:56] ;
assign n305 = LB2D_shift_0[63:56] ;
assign n306 = LB2D_shift_1[63:56] ;
assign n307 = LB2D_shift_2[63:56] ;
assign n308 = LB2D_shift_3[63:56] ;
assign n309 = LB2D_shift_4[63:56] ;
assign n310 = LB2D_shift_5[63:56] ;
assign n311 = LB2D_shift_6[63:56] ;
assign n312 = LB2D_shift_7[63:56] ;
assign n313 =  { ( n311 ) , ( n312 ) }  ;
assign n314 =  { ( n310 ) , ( n313 ) }  ;
assign n315 =  { ( n309 ) , ( n314 ) }  ;
assign n316 =  { ( n308 ) , ( n315 ) }  ;
assign n317 =  { ( n307 ) , ( n316 ) }  ;
assign n318 =  { ( n306 ) , ( n317 ) }  ;
assign n319 =  { ( n305 ) , ( n318 ) }  ;
assign n320 =  { ( n304 ) , ( n319 ) }  ;
assign n321 = n62[55:48] ;
assign n322 = LB2D_shift_0[55:48] ;
assign n323 = LB2D_shift_1[55:48] ;
assign n324 = LB2D_shift_2[55:48] ;
assign n325 = LB2D_shift_3[55:48] ;
assign n326 = LB2D_shift_4[55:48] ;
assign n327 = LB2D_shift_5[55:48] ;
assign n328 = LB2D_shift_6[55:48] ;
assign n329 = LB2D_shift_7[55:48] ;
assign n330 =  { ( n328 ) , ( n329 ) }  ;
assign n331 =  { ( n327 ) , ( n330 ) }  ;
assign n332 =  { ( n326 ) , ( n331 ) }  ;
assign n333 =  { ( n325 ) , ( n332 ) }  ;
assign n334 =  { ( n324 ) , ( n333 ) }  ;
assign n335 =  { ( n323 ) , ( n334 ) }  ;
assign n336 =  { ( n322 ) , ( n335 ) }  ;
assign n337 =  { ( n321 ) , ( n336 ) }  ;
assign n338 = n62[47:40] ;
assign n339 = LB2D_shift_0[47:40] ;
assign n340 = LB2D_shift_1[47:40] ;
assign n341 = LB2D_shift_2[47:40] ;
assign n342 = LB2D_shift_3[47:40] ;
assign n343 = LB2D_shift_4[47:40] ;
assign n344 = LB2D_shift_5[47:40] ;
assign n345 = LB2D_shift_6[47:40] ;
assign n346 = LB2D_shift_7[47:40] ;
assign n347 =  { ( n345 ) , ( n346 ) }  ;
assign n348 =  { ( n344 ) , ( n347 ) }  ;
assign n349 =  { ( n343 ) , ( n348 ) }  ;
assign n350 =  { ( n342 ) , ( n349 ) }  ;
assign n351 =  { ( n341 ) , ( n350 ) }  ;
assign n352 =  { ( n340 ) , ( n351 ) }  ;
assign n353 =  { ( n339 ) , ( n352 ) }  ;
assign n354 =  { ( n338 ) , ( n353 ) }  ;
assign n355 = n62[39:32] ;
assign n356 = LB2D_shift_0[39:32] ;
assign n357 = LB2D_shift_1[39:32] ;
assign n358 = LB2D_shift_2[39:32] ;
assign n359 = LB2D_shift_3[39:32] ;
assign n360 = LB2D_shift_4[39:32] ;
assign n361 = LB2D_shift_5[39:32] ;
assign n362 = LB2D_shift_6[39:32] ;
assign n363 = LB2D_shift_7[39:32] ;
assign n364 =  { ( n362 ) , ( n363 ) }  ;
assign n365 =  { ( n361 ) , ( n364 ) }  ;
assign n366 =  { ( n360 ) , ( n365 ) }  ;
assign n367 =  { ( n359 ) , ( n366 ) }  ;
assign n368 =  { ( n358 ) , ( n367 ) }  ;
assign n369 =  { ( n357 ) , ( n368 ) }  ;
assign n370 =  { ( n356 ) , ( n369 ) }  ;
assign n371 =  { ( n355 ) , ( n370 ) }  ;
assign n372 = n62[31:24] ;
assign n373 = LB2D_shift_0[31:24] ;
assign n374 = LB2D_shift_1[31:24] ;
assign n375 = LB2D_shift_2[31:24] ;
assign n376 = LB2D_shift_3[31:24] ;
assign n377 = LB2D_shift_4[31:24] ;
assign n378 = LB2D_shift_5[31:24] ;
assign n379 = LB2D_shift_6[31:24] ;
assign n380 = LB2D_shift_7[31:24] ;
assign n381 =  { ( n379 ) , ( n380 ) }  ;
assign n382 =  { ( n378 ) , ( n381 ) }  ;
assign n383 =  { ( n377 ) , ( n382 ) }  ;
assign n384 =  { ( n376 ) , ( n383 ) }  ;
assign n385 =  { ( n375 ) , ( n384 ) }  ;
assign n386 =  { ( n374 ) , ( n385 ) }  ;
assign n387 =  { ( n373 ) , ( n386 ) }  ;
assign n388 =  { ( n372 ) , ( n387 ) }  ;
assign n389 = n62[23:16] ;
assign n390 = LB2D_shift_0[23:16] ;
assign n391 = LB2D_shift_1[23:16] ;
assign n392 = LB2D_shift_2[23:16] ;
assign n393 = LB2D_shift_3[23:16] ;
assign n394 = LB2D_shift_4[23:16] ;
assign n395 = LB2D_shift_5[23:16] ;
assign n396 = LB2D_shift_6[23:16] ;
assign n397 = LB2D_shift_7[23:16] ;
assign n398 =  { ( n396 ) , ( n397 ) }  ;
assign n399 =  { ( n395 ) , ( n398 ) }  ;
assign n400 =  { ( n394 ) , ( n399 ) }  ;
assign n401 =  { ( n393 ) , ( n400 ) }  ;
assign n402 =  { ( n392 ) , ( n401 ) }  ;
assign n403 =  { ( n391 ) , ( n402 ) }  ;
assign n404 =  { ( n390 ) , ( n403 ) }  ;
assign n405 =  { ( n389 ) , ( n404 ) }  ;
assign n406 = n62[15:8] ;
assign n407 = LB2D_shift_0[15:8] ;
assign n408 = LB2D_shift_1[15:8] ;
assign n409 = LB2D_shift_2[15:8] ;
assign n410 = LB2D_shift_3[15:8] ;
assign n411 = LB2D_shift_4[15:8] ;
assign n412 = LB2D_shift_5[15:8] ;
assign n413 = LB2D_shift_6[15:8] ;
assign n414 = LB2D_shift_7[15:8] ;
assign n415 =  { ( n413 ) , ( n414 ) }  ;
assign n416 =  { ( n412 ) , ( n415 ) }  ;
assign n417 =  { ( n411 ) , ( n416 ) }  ;
assign n418 =  { ( n410 ) , ( n417 ) }  ;
assign n419 =  { ( n409 ) , ( n418 ) }  ;
assign n420 =  { ( n408 ) , ( n419 ) }  ;
assign n421 =  { ( n407 ) , ( n420 ) }  ;
assign n422 =  { ( n406 ) , ( n421 ) }  ;
assign n423 = n62[7:0] ;
assign n424 = LB2D_shift_0[7:0] ;
assign n425 = LB2D_shift_1[7:0] ;
assign n426 = LB2D_shift_2[7:0] ;
assign n427 = LB2D_shift_3[7:0] ;
assign n428 = LB2D_shift_4[7:0] ;
assign n429 = LB2D_shift_5[7:0] ;
assign n430 = LB2D_shift_6[7:0] ;
assign n431 = LB2D_shift_7[7:0] ;
assign n432 =  { ( n430 ) , ( n431 ) }  ;
assign n433 =  { ( n429 ) , ( n432 ) }  ;
assign n434 =  { ( n428 ) , ( n433 ) }  ;
assign n435 =  { ( n427 ) , ( n434 ) }  ;
assign n436 =  { ( n426 ) , ( n435 ) }  ;
assign n437 =  { ( n425 ) , ( n436 ) }  ;
assign n438 =  { ( n424 ) , ( n437 ) }  ;
assign n439 =  { ( n423 ) , ( n438 ) }  ;
assign n440 =  { ( n422 ) , ( n439 ) }  ;
assign n441 =  { ( n405 ) , ( n440 ) }  ;
assign n442 =  { ( n388 ) , ( n441 ) }  ;
assign n443 =  { ( n371 ) , ( n442 ) }  ;
assign n444 =  { ( n354 ) , ( n443 ) }  ;
assign n445 =  { ( n337 ) , ( n444 ) }  ;
assign n446 =  { ( n320 ) , ( n445 ) }  ;
assign n447 =  { ( n303 ) , ( n446 ) }  ;
assign n448 =  ( n286 ) ? ( n447 ) : ( stencil_stream_buff_0 ) ;
assign n449 =  ( n25 ) ? ( stencil_stream_buff_0 ) : ( stencil_stream_buff_0 ) ;
assign n450 =  ( n22 ) ? ( stencil_stream_buff_0 ) : ( n449 ) ;
assign n451 =  ( n17 ) ? ( n448 ) : ( n450 ) ;
assign n452 =  ( n12 ) ? ( stencil_stream_buff_0 ) : ( n451 ) ;
assign n453 =  ( n9 ) ? ( stencil_stream_buff_0 ) : ( n452 ) ;
assign n454 =  ( n4 ) ? ( stencil_stream_buff_0 ) : ( n453 ) ;
assign n455 =  ( n25 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_1 ) ;
assign n456 =  ( n22 ) ? ( stencil_stream_buff_1 ) : ( n455 ) ;
assign n457 =  ( n17 ) ? ( stencil_stream_buff_0 ) : ( n456 ) ;
assign n458 =  ( n12 ) ? ( stencil_stream_buff_1 ) : ( n457 ) ;
assign n459 =  ( n9 ) ? ( stencil_stream_buff_1 ) : ( n458 ) ;
assign n460 =  ( n4 ) ? ( stencil_stream_buff_1 ) : ( n459 ) ;
assign n461 =  ( n126 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n462 =  ( n15 ) ? ( stencil_stream_empty ) : ( 1'd0 ) ;
assign n463 =  ( n25 ) ? ( stencil_stream_empty ) : ( stencil_stream_empty ) ;
assign n464 =  ( n22 ) ? ( stencil_stream_empty ) : ( n463 ) ;
assign n465 =  ( n17 ) ? ( n462 ) : ( n464 ) ;
assign n466 =  ( n12 ) ? ( n461 ) : ( n465 ) ;
assign n467 =  ( n9 ) ? ( stencil_stream_empty ) : ( n466 ) ;
assign n468 =  ( n4 ) ? ( stencil_stream_empty ) : ( n467 ) ;
assign n469 =  ( stencil_stream_empty ) == ( 1'd1 )  ;
assign n470 =  ( n469 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n471 =  ( n15 ) ? ( stencil_stream_full ) : ( n470 ) ;
assign n472 =  ( n25 ) ? ( stencil_stream_full ) : ( stencil_stream_full ) ;
assign n473 =  ( n22 ) ? ( stencil_stream_full ) : ( n472 ) ;
assign n474 =  ( n17 ) ? ( n471 ) : ( n473 ) ;
assign n475 =  ( n12 ) ? ( 1'd0 ) : ( n474 ) ;
assign n476 =  ( n9 ) ? ( stencil_stream_full ) : ( n475 ) ;
assign n477 =  ( n4 ) ? ( stencil_stream_full ) : ( n476 ) ;
assign n478 = ~ ( n4 ) ;
assign n479 = ~ ( n9 ) ;
assign n480 =  ( n478 ) & ( n479 )  ;
assign n481 = ~ ( n12 ) ;
assign n482 =  ( n480 ) & ( n481 )  ;
assign n483 = ~ ( n17 ) ;
assign n484 =  ( n482 ) & ( n483 )  ;
assign n485 = ~ ( n22 ) ;
assign n486 =  ( n484 ) & ( n485 )  ;
assign n487 = ~ ( n25 ) ;
assign n488 =  ( n486 ) & ( n487 )  ;
assign n489 =  ( n486 ) & ( n25 )  ;
assign n490 =  ( n484 ) & ( n22 )  ;
assign n491 = ~ ( n176 ) ;
assign n492 =  ( n490 ) & ( n491 )  ;
assign n493 =  ( n490 ) & ( n176 )  ;
assign n494 =  ( n482 ) & ( n17 )  ;
assign n495 =  ( n480 ) & ( n12 )  ;
assign n496 =  ( n478 ) & ( n9 )  ;
assign LB2D_proc_0_addr0 = n493 ? (LB2D_proc_x) : (0);
assign LB2D_proc_0_data0 = n493 ? (n175) : (LB2D_proc_0[0]);
assign n497 = ~ ( n178 ) ;
assign n498 =  ( n490 ) & ( n497 )  ;
assign n499 =  ( n490 ) & ( n178 )  ;
assign LB2D_proc_1_addr0 = n499 ? (LB2D_proc_x) : (0);
assign LB2D_proc_1_data0 = n499 ? (n175) : (LB2D_proc_1[0]);
assign n500 = ~ ( n180 ) ;
assign n501 =  ( n490 ) & ( n500 )  ;
assign n502 =  ( n490 ) & ( n180 )  ;
assign LB2D_proc_2_addr0 = n502 ? (LB2D_proc_x) : (0);
assign LB2D_proc_2_data0 = n502 ? (n175) : (LB2D_proc_2[0]);
assign n503 = ~ ( n182 ) ;
assign n504 =  ( n490 ) & ( n503 )  ;
assign n505 =  ( n490 ) & ( n182 )  ;
assign LB2D_proc_3_addr0 = n505 ? (LB2D_proc_x) : (0);
assign LB2D_proc_3_data0 = n505 ? (n175) : (LB2D_proc_3[0]);
assign n506 = ~ ( n184 ) ;
assign n507 =  ( n490 ) & ( n506 )  ;
assign n508 =  ( n490 ) & ( n184 )  ;
assign LB2D_proc_4_addr0 = n508 ? (LB2D_proc_x) : (0);
assign LB2D_proc_4_data0 = n508 ? (n175) : (LB2D_proc_4[0]);
assign n509 = ~ ( n186 ) ;
assign n510 =  ( n490 ) & ( n509 )  ;
assign n511 =  ( n490 ) & ( n186 )  ;
assign LB2D_proc_5_addr0 = n511 ? (LB2D_proc_x) : (0);
assign LB2D_proc_5_data0 = n511 ? (n175) : (LB2D_proc_5[0]);
assign n512 = ~ ( n188 ) ;
assign n513 =  ( n490 ) & ( n512 )  ;
assign n514 =  ( n490 ) & ( n188 )  ;
assign LB2D_proc_6_addr0 = n514 ? (LB2D_proc_x) : (0);
assign LB2D_proc_6_data0 = n514 ? (n175) : (LB2D_proc_6[0]);
assign n515 =  ( LB2D_proc_w ) == ( 64'd7 )  ;
assign n516 = ~ ( n515 ) ;
assign n517 =  ( n490 ) & ( n516 )  ;
assign n518 =  ( n490 ) & ( n515 )  ;
assign LB2D_proc_7_addr0 = n518 ? (LB2D_proc_x) : (0);
assign LB2D_proc_7_data0 = n518 ? (n175) : (LB2D_proc_7[0]);
/*
function [7:0] gb_fun ;
input [647:0] arg0;
    begin
//TODO: Add the specific function HERE.    end
endfunction
*/

always @(posedge clk) begin
   if(rst) begin
       LB1D_buff <= LB1D_buff;
       LB2D_proc_w <= LB2D_proc_w;
       LB2D_proc_x <= LB2D_proc_x;
       LB2D_proc_y <= LB2D_proc_y;
       LB2D_shift_0 <= LB2D_shift_0;
       LB2D_shift_1 <= LB2D_shift_1;
       LB2D_shift_2 <= LB2D_shift_2;
       LB2D_shift_3 <= LB2D_shift_3;
       LB2D_shift_4 <= LB2D_shift_4;
       LB2D_shift_5 <= LB2D_shift_5;
       LB2D_shift_6 <= LB2D_shift_6;
       LB2D_shift_7 <= LB2D_shift_7;
       LB2D_shift_x <= LB2D_shift_x;
       LB2D_shift_y <= LB2D_shift_y;
       arg_0_TDATA <= arg_0_TDATA;
       arg_0_TVALID <= arg_0_TVALID;
       arg_1_TREADY <= arg_1_TREADY;
       in_stream_buff_0 <= in_stream_buff_0;
       in_stream_buff_1 <= in_stream_buff_1;
       in_stream_empty <= in_stream_empty;
       in_stream_full <= in_stream_full;
       slice_stream_buff_0 <= slice_stream_buff_0;
       slice_stream_buff_1 <= slice_stream_buff_1;
       slice_stream_empty <= slice_stream_empty;
       slice_stream_full <= slice_stream_full;
       stencil_stream_buff_0 <= stencil_stream_buff_0;
       stencil_stream_buff_1 <= stencil_stream_buff_1;
       stencil_stream_empty <= stencil_stream_empty;
       stencil_stream_full <= stencil_stream_full;
   end
   else if(step) begin
       LB1D_buff <= n31;
       LB2D_proc_w <= n42;
       LB2D_proc_x <= n50;
       LB2D_proc_y <= n60;
       LB2D_shift_0 <= n68;
       LB2D_shift_1 <= n74;
       LB2D_shift_2 <= n80;
       LB2D_shift_3 <= n86;
       LB2D_shift_4 <= n92;
       LB2D_shift_5 <= n98;
       LB2D_shift_6 <= n104;
       LB2D_shift_7 <= n110;
       LB2D_shift_x <= n119;
       LB2D_shift_y <= n125;
       arg_0_TDATA <= n134;
       arg_0_TVALID <= n140;
       arg_1_TREADY <= n146;
       in_stream_buff_0 <= n152;
       in_stream_buff_1 <= n158;
       in_stream_empty <= n166;
       in_stream_full <= n174;
       slice_stream_buff_0 <= n261;
       slice_stream_buff_1 <= n268;
       slice_stream_empty <= n276;
       slice_stream_full <= n285;
       stencil_stream_buff_0 <= n454;
       stencil_stream_buff_1 <= n460;
       stencil_stream_empty <= n468;
       stencil_stream_full <= n477;
       LB2D_proc_0 [ LB2D_proc_0_addr0 ] <= LB2D_proc_0_data0;
       LB2D_proc_1 [ LB2D_proc_1_addr0 ] <= LB2D_proc_1_data0;
       LB2D_proc_2 [ LB2D_proc_2_addr0 ] <= LB2D_proc_2_data0;
       LB2D_proc_3 [ LB2D_proc_3_addr0 ] <= LB2D_proc_3_data0;
       LB2D_proc_4 [ LB2D_proc_4_addr0 ] <= LB2D_proc_4_data0;
       LB2D_proc_5 [ LB2D_proc_5_addr0 ] <= LB2D_proc_5_data0;
       LB2D_proc_6 [ LB2D_proc_6_addr0 ] <= LB2D_proc_6_data0;
       LB2D_proc_7 [ LB2D_proc_7_addr0 ] <= LB2D_proc_7_data0;
   end
end
endmodule
