module SPEC_B(
arg_0_TREADY,
arg_1_TDATA,
arg_1_TVALID,
LB1D_buff,
LB1D_in,
LB1D_it_1,
LB1D_p_cnt,
LB1D_uIn,
LB2D_proc_w,
LB2D_proc_x,
LB2D_proc_y,
LB2D_shift_0,
LB2D_shift_1,
LB2D_shift_2,
LB2D_shift_3,
LB2D_shift_4,
LB2D_shift_5,
LB2D_shift_6,
LB2D_shift_7,
LB2D_shift_x,
LB2D_shift_y,
arg_0_TDATA,
arg_0_TVALID,
arg_1_TREADY,
gb_exit_it_1,
gb_exit_it_2,
gb_exit_it_3,
gb_exit_it_4,
gb_exit_it_5,
gb_exit_it_6,
gb_exit_it_7,
gb_exit_it_8,
gb_p_cnt,
gb_pp_it_1,
gb_pp_it_2,
gb_pp_it_3,
gb_pp_it_4,
gb_pp_it_5,
gb_pp_it_6,
gb_pp_it_7,
gb_pp_it_8,
gb_pp_it_9,
in_stream_buff_0,
in_stream_buff_1,
in_stream_empty,
in_stream_full,
slice_stream_buff_0,
slice_stream_buff_1,
slice_stream_empty,
slice_stream_full,
stencil_stream_buff_0,
stencil_stream_buff_1,
stencil_stream_empty,
stencil_stream_full,
clk,rst,
step
);
input            arg_0_TREADY;
input      [7:0] arg_1_TDATA;
input            arg_1_TVALID;
input clk;
input rst;
input step;
output      [7:0] LB1D_buff;
output      [7:0] LB1D_in;
output            LB1D_it_1;
output     [18:0] LB1D_p_cnt;
output      [7:0] LB1D_uIn;
output     [63:0] LB2D_proc_w;
output      [8:0] LB2D_proc_x;
output      [9:0] LB2D_proc_y;
output     [71:0] LB2D_shift_0;
output     [71:0] LB2D_shift_1;
output     [71:0] LB2D_shift_2;
output     [71:0] LB2D_shift_3;
output     [71:0] LB2D_shift_4;
output     [71:0] LB2D_shift_5;
output     [71:0] LB2D_shift_6;
output     [71:0] LB2D_shift_7;
output      [8:0] LB2D_shift_x;
output      [9:0] LB2D_shift_y;
output      [7:0] arg_0_TDATA;
output            arg_0_TVALID;
output            arg_1_TREADY;
output            gb_exit_it_1;
output            gb_exit_it_2;
output            gb_exit_it_3;
output            gb_exit_it_4;
output            gb_exit_it_5;
output            gb_exit_it_6;
output            gb_exit_it_7;
output            gb_exit_it_8;
output     [18:0] gb_p_cnt;
output            gb_pp_it_1;
output            gb_pp_it_2;
output            gb_pp_it_3;
output            gb_pp_it_4;
output            gb_pp_it_5;
output            gb_pp_it_6;
output            gb_pp_it_7;
output            gb_pp_it_8;
output            gb_pp_it_9;
output      [7:0] in_stream_buff_0;
output      [7:0] in_stream_buff_1;
output            in_stream_empty;
output            in_stream_full;
output     [71:0] slice_stream_buff_0;
output     [71:0] slice_stream_buff_1;
output            slice_stream_empty;
output            slice_stream_full;
output    [647:0] stencil_stream_buff_0;
output    [647:0] stencil_stream_buff_1;
output            stencil_stream_empty;
output            stencil_stream_full;
reg      [7:0] LB1D_buff;
reg      [7:0] LB1D_in;
reg            LB1D_it_1;
reg     [18:0] LB1D_p_cnt;
reg      [7:0] LB1D_uIn;
reg     [63:0] LB2D_proc_w;
reg      [8:0] LB2D_proc_x;
reg      [9:0] LB2D_proc_y;
reg     [71:0] LB2D_shift_0;
reg     [71:0] LB2D_shift_1;
reg     [71:0] LB2D_shift_2;
reg     [71:0] LB2D_shift_3;
reg     [71:0] LB2D_shift_4;
reg     [71:0] LB2D_shift_5;
reg     [71:0] LB2D_shift_6;
reg     [71:0] LB2D_shift_7;
reg      [8:0] LB2D_shift_x;
reg      [9:0] LB2D_shift_y;
reg      [7:0] arg_0_TDATA;
reg            arg_0_TVALID;
reg            arg_1_TREADY;
reg            gb_exit_it_1;
reg            gb_exit_it_2;
reg            gb_exit_it_3;
reg            gb_exit_it_4;
reg            gb_exit_it_5;
reg            gb_exit_it_6;
reg            gb_exit_it_7;
reg            gb_exit_it_8;
reg     [18:0] gb_p_cnt;
reg            gb_pp_it_1;
reg            gb_pp_it_2;
reg            gb_pp_it_3;
reg            gb_pp_it_4;
reg            gb_pp_it_5;
reg            gb_pp_it_6;
reg            gb_pp_it_7;
reg            gb_pp_it_8;
reg            gb_pp_it_9;
reg      [7:0] in_stream_buff_0;
reg      [7:0] in_stream_buff_1;
reg            in_stream_empty;
reg            in_stream_full;
reg     [71:0] slice_stream_buff_0;
reg     [71:0] slice_stream_buff_1;
reg            slice_stream_empty;
reg            slice_stream_full;
reg    [647:0] stencil_stream_buff_0;
reg    [647:0] stencil_stream_buff_1;
reg            stencil_stream_empty;
reg            stencil_stream_full;
wire            arg_0_TREADY;
wire      [7:0] arg_1_TDATA;
wire            arg_1_TVALID;
wire            n0;
wire            n1;
wire            n2;
wire            n3;
wire            n4;
wire            n5;
wire            n6;
wire            n7;
wire            n8;
wire            n9;
wire            n10;
wire            n11;
wire            n12;
wire            n13;
wire            n14;
wire            n15;
wire            n16;
wire            n17;
wire            n18;
wire            n19;
wire            n20;
wire            n21;
wire            n22;
wire            n23;
wire            n24;
wire            n25;
wire            n26;
wire            n27;
wire            n28;
wire            n29;
wire            n30;
wire            n31;
wire            n32;
wire            n33;
wire            n34;
wire            n35;
wire            n36;
wire            n37;
wire            n38;
wire            n39;
wire      [7:0] n40;
wire      [7:0] n41;
wire      [7:0] n42;
wire      [7:0] n43;
wire      [7:0] n44;
wire      [7:0] n45;
wire      [7:0] n46;
wire      [7:0] n47;
wire      [7:0] n48;
wire      [7:0] n49;
wire      [7:0] n50;
wire      [7:0] n51;
wire      [7:0] n52;
wire      [7:0] n53;
wire            n54;
wire            n55;
wire            n56;
wire     [18:0] n57;
wire     [18:0] n58;
wire     [18:0] n59;
wire     [18:0] n60;
wire     [18:0] n61;
wire     [18:0] n62;
wire     [18:0] n63;
wire     [18:0] n64;
wire      [7:0] n65;
wire      [7:0] n66;
wire      [7:0] n67;
wire      [7:0] n68;
wire      [7:0] n69;
wire      [7:0] n70;
wire            n71;
wire            n72;
wire     [63:0] n73;
wire     [63:0] n74;
wire     [63:0] n75;
wire     [63:0] n76;
wire     [63:0] n77;
wire     [63:0] n78;
wire     [63:0] n79;
wire     [63:0] n80;
wire     [63:0] n81;
wire      [8:0] n82;
wire      [8:0] n83;
wire      [8:0] n84;
wire      [8:0] n85;
wire      [8:0] n86;
wire      [8:0] n87;
wire      [8:0] n88;
wire      [8:0] n89;
wire            n90;
wire      [9:0] n91;
wire      [9:0] n92;
wire      [9:0] n93;
wire      [9:0] n94;
wire      [9:0] n95;
wire      [9:0] n96;
wire      [9:0] n97;
wire      [9:0] n98;
wire      [9:0] n99;
wire     [71:0] n100;
wire     [71:0] n101;
wire     [71:0] n102;
wire     [71:0] n103;
wire     [71:0] n104;
wire     [71:0] n105;
wire     [71:0] n106;
wire     [71:0] n107;
wire     [71:0] n108;
wire     [71:0] n109;
wire     [71:0] n110;
wire     [71:0] n111;
wire     [71:0] n112;
wire     [71:0] n113;
wire     [71:0] n114;
wire     [71:0] n115;
wire     [71:0] n116;
wire     [71:0] n117;
wire     [71:0] n118;
wire     [71:0] n119;
wire     [71:0] n120;
wire     [71:0] n121;
wire     [71:0] n122;
wire     [71:0] n123;
wire     [71:0] n124;
wire     [71:0] n125;
wire     [71:0] n126;
wire     [71:0] n127;
wire     [71:0] n128;
wire     [71:0] n129;
wire     [71:0] n130;
wire     [71:0] n131;
wire     [71:0] n132;
wire     [71:0] n133;
wire     [71:0] n134;
wire     [71:0] n135;
wire     [71:0] n136;
wire     [71:0] n137;
wire     [71:0] n138;
wire     [71:0] n139;
wire     [71:0] n140;
wire     [71:0] n141;
wire            n142;
wire     [71:0] n143;
wire     [71:0] n144;
wire     [71:0] n145;
wire     [71:0] n146;
wire     [71:0] n147;
wire     [71:0] n148;
wire     [71:0] n149;
wire            n150;
wire            n151;
wire            n152;
wire            n153;
wire      [8:0] n154;
wire      [8:0] n155;
wire      [8:0] n156;
wire      [8:0] n157;
wire      [8:0] n158;
wire      [8:0] n159;
wire      [8:0] n160;
wire      [8:0] n161;
wire            n162;
wire            n163;
wire      [9:0] n164;
wire      [9:0] n165;
wire      [9:0] n166;
wire      [9:0] n167;
wire      [9:0] n168;
wire      [9:0] n169;
wire      [9:0] n170;
wire      [9:0] n171;
wire      [9:0] n172;
wire            n173;
wire    [647:0] n174;
wire      [7:0] n175;
wire      [7:0] n176;
wire      [7:0] n177;
wire      [7:0] n178;
wire      [7:0] n179;
wire      [7:0] n180;
wire      [7:0] n181;
wire            n182;
wire            n183;
wire            n184;
wire            n185;
wire            n186;
wire            n187;
wire            n188;
wire            n189;
wire            n190;
wire            n191;
wire            n192;
wire            n193;
wire            n194;
wire            n195;
wire            n196;
wire            n197;
wire            n198;
wire            n199;
wire            n200;
wire            n201;
wire            n202;
wire            n203;
wire            n204;
wire            n205;
wire            n206;
wire            n207;
wire            n208;
wire            n209;
wire            n210;
wire            n211;
wire            n212;
wire            n213;
wire            n214;
wire            n215;
wire            n216;
wire            n217;
wire            n218;
wire            n219;
wire            n220;
wire            n221;
wire            n222;
wire            n223;
wire            n224;
wire            n225;
wire            n226;
wire            n227;
wire            n228;
wire            n229;
wire            n230;
wire            n231;
wire            n232;
wire            n233;
wire            n234;
wire            n235;
wire            n236;
wire            n237;
wire            n238;
wire            n239;
wire            n240;
wire            n241;
wire            n242;
wire            n243;
wire            n244;
wire            n245;
wire            n246;
wire            n247;
wire     [18:0] n248;
wire     [18:0] n249;
wire     [18:0] n250;
wire     [18:0] n251;
wire     [18:0] n252;
wire     [18:0] n253;
wire     [18:0] n254;
wire     [18:0] n255;
wire            n256;
wire            n257;
wire            n258;
wire            n259;
wire            n260;
wire            n261;
wire            n262;
wire            n263;
wire            n264;
wire            n265;
wire            n266;
wire            n267;
wire            n268;
wire            n269;
wire            n270;
wire            n271;
wire            n272;
wire            n273;
wire            n274;
wire            n275;
wire            n276;
wire            n277;
wire            n278;
wire            n279;
wire            n280;
wire            n281;
wire            n282;
wire            n283;
wire            n284;
wire            n285;
wire            n286;
wire            n287;
wire            n288;
wire            n289;
wire            n290;
wire            n291;
wire            n292;
wire            n293;
wire            n294;
wire            n295;
wire            n296;
wire            n297;
wire            n298;
wire            n299;
wire            n300;
wire            n301;
wire            n302;
wire            n303;
wire            n304;
wire            n305;
wire            n306;
wire            n307;
wire            n308;
wire            n309;
wire      [7:0] n310;
wire      [7:0] n311;
wire      [7:0] n312;
wire      [7:0] n313;
wire      [7:0] n314;
wire      [7:0] n315;
wire      [7:0] n316;
wire      [7:0] n317;
wire      [7:0] n318;
wire      [7:0] n319;
wire      [7:0] n320;
wire      [7:0] n321;
wire            n322;
wire            n323;
wire            n324;
wire            n325;
wire            n326;
wire            n327;
wire            n328;
wire            n329;
wire            n330;
wire            n331;
wire            n332;
wire            n333;
wire            n334;
wire            n335;
wire            n336;
wire            n337;
wire      [7:0] n338;
wire            n339;
wire      [8:0] n340;
wire      [7:0] n341;
wire            n342;
wire      [7:0] n343;
wire            n344;
wire      [7:0] n345;
wire            n346;
wire      [7:0] n347;
wire            n348;
wire      [7:0] n349;
wire            n350;
wire      [7:0] n351;
wire            n352;
wire      [7:0] n353;
wire      [7:0] n354;
wire      [7:0] n355;
wire      [7:0] n356;
wire      [7:0] n357;
wire      [7:0] n358;
wire      [7:0] n359;
wire      [7:0] n360;
wire      [7:0] n361;
wire      [7:0] n362;
wire      [7:0] n363;
wire      [7:0] n364;
wire      [7:0] n365;
wire      [7:0] n366;
wire      [7:0] n367;
wire      [7:0] n368;
wire      [7:0] n369;
wire      [7:0] n370;
wire      [7:0] n371;
wire      [7:0] n372;
wire      [7:0] n373;
wire      [7:0] n374;
wire      [7:0] n375;
wire      [7:0] n376;
wire      [7:0] n377;
wire      [7:0] n378;
wire      [7:0] n379;
wire      [7:0] n380;
wire      [7:0] n381;
wire      [7:0] n382;
wire      [7:0] n383;
wire      [7:0] n384;
wire      [7:0] n385;
wire      [7:0] n386;
wire      [7:0] n387;
wire      [7:0] n388;
wire      [7:0] n389;
wire      [7:0] n390;
wire      [7:0] n391;
wire      [7:0] n392;
wire      [7:0] n393;
wire      [7:0] n394;
wire      [7:0] n395;
wire      [7:0] n396;
wire      [7:0] n397;
wire      [7:0] n398;
wire      [7:0] n399;
wire      [7:0] n400;
wire      [7:0] n401;
wire      [7:0] n402;
wire      [7:0] n403;
wire      [7:0] n404;
wire      [7:0] n405;
wire      [7:0] n406;
wire      [7:0] n407;
wire      [7:0] n408;
wire      [7:0] n409;
wire      [7:0] n410;
wire     [15:0] n411;
wire     [23:0] n412;
wire     [31:0] n413;
wire     [39:0] n414;
wire     [47:0] n415;
wire     [55:0] n416;
wire     [63:0] n417;
wire     [71:0] n418;
wire     [71:0] n419;
wire     [71:0] n420;
wire     [71:0] n421;
wire     [71:0] n422;
wire     [71:0] n423;
wire     [71:0] n424;
wire     [71:0] n425;
wire     [71:0] n426;
wire     [71:0] n427;
wire     [71:0] n428;
wire     [71:0] n429;
wire     [71:0] n430;
wire     [71:0] n431;
wire     [71:0] n432;
wire            n433;
wire            n434;
wire            n435;
wire            n436;
wire            n437;
wire            n438;
wire            n439;
wire            n440;
wire            n441;
wire            n442;
wire            n443;
wire            n444;
wire            n445;
wire            n446;
wire            n447;
wire            n448;
wire            n449;
wire            n450;
wire            n451;
wire            n452;
wire      [7:0] n453;
wire      [7:0] n454;
wire      [7:0] n455;
wire      [7:0] n456;
wire      [7:0] n457;
wire      [7:0] n458;
wire      [7:0] n459;
wire      [7:0] n460;
wire      [7:0] n461;
wire     [15:0] n462;
wire     [23:0] n463;
wire     [31:0] n464;
wire     [39:0] n465;
wire     [47:0] n466;
wire     [55:0] n467;
wire     [63:0] n468;
wire     [71:0] n469;
wire      [7:0] n470;
wire      [7:0] n471;
wire      [7:0] n472;
wire      [7:0] n473;
wire      [7:0] n474;
wire      [7:0] n475;
wire      [7:0] n476;
wire      [7:0] n477;
wire      [7:0] n478;
wire     [15:0] n479;
wire     [23:0] n480;
wire     [31:0] n481;
wire     [39:0] n482;
wire     [47:0] n483;
wire     [55:0] n484;
wire     [63:0] n485;
wire     [71:0] n486;
wire      [7:0] n487;
wire      [7:0] n488;
wire      [7:0] n489;
wire      [7:0] n490;
wire      [7:0] n491;
wire      [7:0] n492;
wire      [7:0] n493;
wire      [7:0] n494;
wire      [7:0] n495;
wire     [15:0] n496;
wire     [23:0] n497;
wire     [31:0] n498;
wire     [39:0] n499;
wire     [47:0] n500;
wire     [55:0] n501;
wire     [63:0] n502;
wire     [71:0] n503;
wire      [7:0] n504;
wire      [7:0] n505;
wire      [7:0] n506;
wire      [7:0] n507;
wire      [7:0] n508;
wire      [7:0] n509;
wire      [7:0] n510;
wire      [7:0] n511;
wire      [7:0] n512;
wire     [15:0] n513;
wire     [23:0] n514;
wire     [31:0] n515;
wire     [39:0] n516;
wire     [47:0] n517;
wire     [55:0] n518;
wire     [63:0] n519;
wire     [71:0] n520;
wire      [7:0] n521;
wire      [7:0] n522;
wire      [7:0] n523;
wire      [7:0] n524;
wire      [7:0] n525;
wire      [7:0] n526;
wire      [7:0] n527;
wire      [7:0] n528;
wire      [7:0] n529;
wire     [15:0] n530;
wire     [23:0] n531;
wire     [31:0] n532;
wire     [39:0] n533;
wire     [47:0] n534;
wire     [55:0] n535;
wire     [63:0] n536;
wire     [71:0] n537;
wire      [7:0] n538;
wire      [7:0] n539;
wire      [7:0] n540;
wire      [7:0] n541;
wire      [7:0] n542;
wire      [7:0] n543;
wire      [7:0] n544;
wire      [7:0] n545;
wire      [7:0] n546;
wire     [15:0] n547;
wire     [23:0] n548;
wire     [31:0] n549;
wire     [39:0] n550;
wire     [47:0] n551;
wire     [55:0] n552;
wire     [63:0] n553;
wire     [71:0] n554;
wire      [7:0] n555;
wire      [7:0] n556;
wire      [7:0] n557;
wire      [7:0] n558;
wire      [7:0] n559;
wire      [7:0] n560;
wire      [7:0] n561;
wire      [7:0] n562;
wire      [7:0] n563;
wire     [15:0] n564;
wire     [23:0] n565;
wire     [31:0] n566;
wire     [39:0] n567;
wire     [47:0] n568;
wire     [55:0] n569;
wire     [63:0] n570;
wire     [71:0] n571;
wire      [7:0] n572;
wire      [7:0] n573;
wire      [7:0] n574;
wire      [7:0] n575;
wire      [7:0] n576;
wire      [7:0] n577;
wire      [7:0] n578;
wire      [7:0] n579;
wire      [7:0] n580;
wire     [15:0] n581;
wire     [23:0] n582;
wire     [31:0] n583;
wire     [39:0] n584;
wire     [47:0] n585;
wire     [55:0] n586;
wire     [63:0] n587;
wire     [71:0] n588;
wire      [7:0] n589;
wire      [7:0] n590;
wire      [7:0] n591;
wire      [7:0] n592;
wire      [7:0] n593;
wire      [7:0] n594;
wire      [7:0] n595;
wire      [7:0] n596;
wire      [7:0] n597;
wire     [15:0] n598;
wire     [23:0] n599;
wire     [31:0] n600;
wire     [39:0] n601;
wire     [47:0] n602;
wire     [55:0] n603;
wire     [63:0] n604;
wire     [71:0] n605;
wire    [143:0] n606;
wire    [215:0] n607;
wire    [287:0] n608;
wire    [359:0] n609;
wire    [431:0] n610;
wire    [503:0] n611;
wire    [575:0] n612;
wire    [647:0] n613;
wire    [647:0] n614;
wire    [647:0] n615;
wire    [647:0] n616;
wire    [647:0] n617;
wire    [647:0] n618;
wire    [647:0] n619;
wire    [647:0] n620;
wire    [647:0] n621;
wire    [647:0] n622;
wire    [647:0] n623;
wire    [647:0] n624;
wire    [647:0] n625;
wire    [647:0] n626;
wire            n627;
wire            n628;
wire            n629;
wire            n630;
wire            n631;
wire            n632;
wire            n633;
wire            n634;
wire            n635;
wire            n636;
wire            n637;
wire            n638;
wire            n639;
wire            n640;
wire            n641;
wire            n642;
wire            n643;
wire            n644;
wire            n645;
wire      [8:0] LB2D_proc_0_addr0;
wire      [7:0] LB2D_proc_0_data0;
wire            n646;
wire            n647;
wire            n648;
wire            n649;
wire            n650;
wire            n651;
wire            n652;
wire            n653;
wire            n654;
wire            n655;
wire            n656;
wire            n657;
wire            n658;
wire            n659;
wire            n660;
wire            n661;
wire            n662;
wire            n663;
wire            n664;
wire      [8:0] LB2D_proc_1_addr0;
wire      [7:0] LB2D_proc_1_data0;
wire            n665;
wire            n666;
wire            n667;
wire      [8:0] LB2D_proc_2_addr0;
wire      [7:0] LB2D_proc_2_data0;
wire            n668;
wire            n669;
wire            n670;
wire      [8:0] LB2D_proc_3_addr0;
wire      [7:0] LB2D_proc_3_data0;
wire            n671;
wire            n672;
wire            n673;
wire      [8:0] LB2D_proc_4_addr0;
wire      [7:0] LB2D_proc_4_data0;
wire            n674;
wire            n675;
wire            n676;
wire      [8:0] LB2D_proc_5_addr0;
wire      [7:0] LB2D_proc_5_data0;
wire            n677;
wire            n678;
wire            n679;
wire      [8:0] LB2D_proc_6_addr0;
wire      [7:0] LB2D_proc_6_data0;
wire            n680;
wire            n681;
wire            n682;
wire      [8:0] LB2D_proc_7_addr0;
wire      [7:0] LB2D_proc_7_data0;
wire            n683;
wire            n684;
wire            n685;
reg      [7:0] LB2D_proc_0[511:0];
reg      [7:0] LB2D_proc_1[511:0];
reg      [7:0] LB2D_proc_2[511:0];
reg      [7:0] LB2D_proc_3[511:0];
reg      [7:0] LB2D_proc_4[511:0];
reg      [7:0] LB2D_proc_5[511:0];
reg      [7:0] LB2D_proc_6[511:0];
reg      [7:0] LB2D_proc_7[511:0];
wire clk;
wire rst;
wire step;
assign n0 =  ( arg_1_TREADY ) == ( 1'd1 )  ;
assign n1 =  ( in_stream_full ) == ( 1'd0 )  ;
assign n2 =  ( n0 ) & ( n1 )  ;
assign n3 =  ( LB1D_it_1 ) == ( 1'd1 )  ;
assign n4 =  ( n2 ) & ( n3 )  ;
assign n5 =  ( LB1D_p_cnt ) == ( 19'd316224 )  ;
assign n6 =  ( n4 ) & ( n5 )  ;
assign n7 =  ( arg_0_TREADY ) == ( 1'd1 )  ;
assign n8 =  ( arg_0_TVALID ) == ( 1'd1 )  ;
assign n9 =  ( n7 ) & ( n8 )  ;
assign n10 =  ( arg_1_TVALID ) == ( 1'd0 )  ;
assign n11 =  ( n9 ) & ( n10 )  ;
assign n12 =  ( arg_0_TVALID ) == ( 1'd0 )  ;
assign n13 =  ( gb_exit_it_1 ) == ( 1'd0 )  ;
assign n14 =  ( stencil_stream_empty ) == ( 1'd0 )  ;
assign n15 =  ( n13 ) & ( n14 )  ;
assign n16 =  ( gb_exit_it_1 ) == ( 1'd1 )  ;
assign n17 =  ( gb_exit_it_8 ) == ( 1'd0 )  ;
assign n18 =  ( n16 ) & ( n17 )  ;
assign n19 =  ( n15 ) | ( n18 )  ;
assign n20 =  ( n12 ) & ( n19 )  ;
assign n21 =  ( slice_stream_empty ) == ( 1'd0 )  ;
assign n22 =  ( LB2D_shift_x ) != ( 9'd488 )  ;
assign n23 =  ( n21 ) & ( n22 )  ;
assign n24 =  ( stencil_stream_full ) == ( 1'd0 )  ;
assign n25 =  ( LB2D_shift_x ) < ( 9'd8 )  ;
assign n26 =  ( LB2D_shift_x ) > ( 9'd0 )  ;
assign n27 =  ( n25 ) & ( n26 )  ;
assign n28 =  ( n24 ) | ( n27 )  ;
assign n29 =  ( n23 ) & ( n28 )  ;
assign n30 =  ( in_stream_empty ) == ( 1'd0 )  ;
assign n31 =  ( slice_stream_full ) == ( 1'd0 )  ;
assign n32 =  ( LB2D_proc_y ) < ( 10'd8 )  ;
assign n33 =  ( n31 ) | ( n32 )  ;
assign n34 =  ( n30 ) & ( n33 )  ;
assign n35 =  ( arg_1_TREADY ) == ( 1'd0 )  ;
assign n36 =  ( n35 ) & ( n1 )  ;
assign n37 =  ( LB1D_it_1 ) == ( 1'd0 )  ;
assign n38 =  ( n36 ) & ( n37 )  ;
assign n39 =  ( n36 ) & ( n3 )  ;
assign n40 =  ( n39 ) ? ( LB1D_uIn ) : ( LB1D_buff ) ;
assign n41 =  ( n38 ) ? ( LB1D_uIn ) : ( n40 ) ;
assign n42 =  ( n34 ) ? ( LB1D_buff ) : ( n41 ) ;
assign n43 =  ( n29 ) ? ( LB1D_buff ) : ( n42 ) ;
assign n44 =  ( n20 ) ? ( LB1D_buff ) : ( n43 ) ;
assign n45 =  ( n11 ) ? ( LB1D_buff ) : ( n44 ) ;
assign n46 =  ( n6 ) ? ( LB1D_uIn ) : ( n45 ) ;
assign n47 =  ( n39 ) ? ( LB1D_in ) : ( LB1D_in ) ;
assign n48 =  ( n38 ) ? ( LB1D_in ) : ( n47 ) ;
assign n49 =  ( n34 ) ? ( LB1D_in ) : ( n48 ) ;
assign n50 =  ( n29 ) ? ( LB1D_in ) : ( n49 ) ;
assign n51 =  ( n20 ) ? ( LB1D_in ) : ( n50 ) ;
assign n52 =  ( n11 ) ? ( LB1D_in ) : ( n51 ) ;
assign n53 =  ( n6 ) ? ( LB1D_in ) : ( n52 ) ;
assign n54 =  ( n39 ) ? ( 1'd1 ) : ( LB1D_it_1 ) ;
assign n55 =  ( n38 ) ? ( 1'd1 ) : ( n54 ) ;
assign n56 =  ( n6 ) ? ( 1'd0 ) : ( n55 ) ;
assign n57 =  ( LB1D_p_cnt ) + ( 19'd1 )  ;
assign n58 =  ( n39 ) ? ( n57 ) : ( LB1D_p_cnt ) ;
assign n59 =  ( n38 ) ? ( n57 ) : ( n58 ) ;
assign n60 =  ( n34 ) ? ( LB1D_p_cnt ) : ( n59 ) ;
assign n61 =  ( n29 ) ? ( LB1D_p_cnt ) : ( n60 ) ;
assign n62 =  ( n20 ) ? ( LB1D_p_cnt ) : ( n61 ) ;
assign n63 =  ( n11 ) ? ( LB1D_p_cnt ) : ( n62 ) ;
assign n64 =  ( n6 ) ? ( 19'd0 ) : ( n63 ) ;
assign n65 =  ( n39 ) ? ( LB1D_in ) : ( LB1D_uIn ) ;
assign n66 =  ( n38 ) ? ( LB1D_in ) : ( n65 ) ;
assign n67 =  ( n34 ) ? ( LB1D_uIn ) : ( n66 ) ;
assign n68 =  ( n29 ) ? ( LB1D_uIn ) : ( n67 ) ;
assign n69 =  ( n20 ) ? ( LB1D_uIn ) : ( n68 ) ;
assign n70 =  ( n6 ) ? ( LB1D_in ) : ( n69 ) ;
assign n71 =  ( LB2D_proc_x ) == ( 9'd488 )  ;
assign n72 =  ( LB2D_proc_w ) == ( 64'd7 )  ;
assign n73 =  ( LB2D_proc_w ) + ( 64'd1 )  ;
assign n74 =  ( n72 ) ? ( 64'd0 ) : ( n73 ) ;
assign n75 =  ( n71 ) ? ( n74 ) : ( LB2D_proc_w ) ;
assign n76 =  ( n39 ) ? ( LB2D_proc_w ) : ( LB2D_proc_w ) ;
assign n77 =  ( n34 ) ? ( n75 ) : ( n76 ) ;
assign n78 =  ( n29 ) ? ( LB2D_proc_w ) : ( n77 ) ;
assign n79 =  ( n20 ) ? ( LB2D_proc_w ) : ( n78 ) ;
assign n80 =  ( n11 ) ? ( LB2D_proc_w ) : ( n79 ) ;
assign n81 =  ( n6 ) ? ( LB2D_proc_w ) : ( n80 ) ;
assign n82 =  ( LB2D_proc_x ) + ( 9'd1 )  ;
assign n83 =  ( n71 ) ? ( 9'd1 ) : ( n82 ) ;
assign n84 =  ( n39 ) ? ( LB2D_proc_x ) : ( LB2D_proc_x ) ;
assign n85 =  ( n34 ) ? ( n83 ) : ( n84 ) ;
assign n86 =  ( n29 ) ? ( LB2D_proc_x ) : ( n85 ) ;
assign n87 =  ( n20 ) ? ( LB2D_proc_x ) : ( n86 ) ;
assign n88 =  ( n11 ) ? ( LB2D_proc_x ) : ( n87 ) ;
assign n89 =  ( n6 ) ? ( LB2D_proc_x ) : ( n88 ) ;
assign n90 =  ( LB2D_proc_y ) == ( 10'd648 )  ;
assign n91 =  ( LB2D_proc_y ) + ( 10'd1 )  ;
assign n92 =  ( n90 ) ? ( 10'd0 ) : ( n91 ) ;
assign n93 =  ( n71 ) ? ( n92 ) : ( LB2D_proc_y ) ;
assign n94 =  ( n39 ) ? ( LB2D_proc_y ) : ( LB2D_proc_y ) ;
assign n95 =  ( n34 ) ? ( n93 ) : ( n94 ) ;
assign n96 =  ( n29 ) ? ( LB2D_proc_y ) : ( n95 ) ;
assign n97 =  ( n20 ) ? ( LB2D_proc_y ) : ( n96 ) ;
assign n98 =  ( n11 ) ? ( LB2D_proc_y ) : ( n97 ) ;
assign n99 =  ( n6 ) ? ( LB2D_proc_y ) : ( n98 ) ;
assign n100 =  ( n39 ) ? ( LB2D_shift_0 ) : ( LB2D_shift_0 ) ;
assign n101 =  ( n34 ) ? ( LB2D_shift_0 ) : ( n100 ) ;
assign n102 =  ( n29 ) ? ( LB2D_shift_1 ) : ( n101 ) ;
assign n103 =  ( n20 ) ? ( LB2D_shift_0 ) : ( n102 ) ;
assign n104 =  ( n11 ) ? ( LB2D_shift_0 ) : ( n103 ) ;
assign n105 =  ( n6 ) ? ( LB2D_shift_0 ) : ( n104 ) ;
assign n106 =  ( n39 ) ? ( LB2D_shift_1 ) : ( LB2D_shift_1 ) ;
assign n107 =  ( n34 ) ? ( LB2D_shift_1 ) : ( n106 ) ;
assign n108 =  ( n29 ) ? ( LB2D_shift_2 ) : ( n107 ) ;
assign n109 =  ( n20 ) ? ( LB2D_shift_1 ) : ( n108 ) ;
assign n110 =  ( n11 ) ? ( LB2D_shift_1 ) : ( n109 ) ;
assign n111 =  ( n6 ) ? ( LB2D_shift_1 ) : ( n110 ) ;
assign n112 =  ( n39 ) ? ( LB2D_shift_2 ) : ( LB2D_shift_2 ) ;
assign n113 =  ( n34 ) ? ( LB2D_shift_2 ) : ( n112 ) ;
assign n114 =  ( n29 ) ? ( LB2D_shift_3 ) : ( n113 ) ;
assign n115 =  ( n20 ) ? ( LB2D_shift_2 ) : ( n114 ) ;
assign n116 =  ( n11 ) ? ( LB2D_shift_2 ) : ( n115 ) ;
assign n117 =  ( n6 ) ? ( LB2D_shift_2 ) : ( n116 ) ;
assign n118 =  ( n39 ) ? ( LB2D_shift_3 ) : ( LB2D_shift_3 ) ;
assign n119 =  ( n34 ) ? ( LB2D_shift_3 ) : ( n118 ) ;
assign n120 =  ( n29 ) ? ( LB2D_shift_4 ) : ( n119 ) ;
assign n121 =  ( n20 ) ? ( LB2D_shift_3 ) : ( n120 ) ;
assign n122 =  ( n11 ) ? ( LB2D_shift_3 ) : ( n121 ) ;
assign n123 =  ( n6 ) ? ( LB2D_shift_3 ) : ( n122 ) ;
assign n124 =  ( n39 ) ? ( LB2D_shift_4 ) : ( LB2D_shift_4 ) ;
assign n125 =  ( n34 ) ? ( LB2D_shift_4 ) : ( n124 ) ;
assign n126 =  ( n29 ) ? ( LB2D_shift_5 ) : ( n125 ) ;
assign n127 =  ( n20 ) ? ( LB2D_shift_4 ) : ( n126 ) ;
assign n128 =  ( n11 ) ? ( LB2D_shift_4 ) : ( n127 ) ;
assign n129 =  ( n6 ) ? ( LB2D_shift_4 ) : ( n128 ) ;
assign n130 =  ( n39 ) ? ( LB2D_shift_5 ) : ( LB2D_shift_5 ) ;
assign n131 =  ( n34 ) ? ( LB2D_shift_5 ) : ( n130 ) ;
assign n132 =  ( n29 ) ? ( LB2D_shift_6 ) : ( n131 ) ;
assign n133 =  ( n20 ) ? ( LB2D_shift_5 ) : ( n132 ) ;
assign n134 =  ( n11 ) ? ( LB2D_shift_5 ) : ( n133 ) ;
assign n135 =  ( n6 ) ? ( LB2D_shift_5 ) : ( n134 ) ;
assign n136 =  ( n39 ) ? ( LB2D_shift_6 ) : ( LB2D_shift_6 ) ;
assign n137 =  ( n34 ) ? ( LB2D_shift_6 ) : ( n136 ) ;
assign n138 =  ( n29 ) ? ( LB2D_shift_7 ) : ( n137 ) ;
assign n139 =  ( n20 ) ? ( LB2D_shift_6 ) : ( n138 ) ;
assign n140 =  ( n11 ) ? ( LB2D_shift_6 ) : ( n139 ) ;
assign n141 =  ( n6 ) ? ( LB2D_shift_6 ) : ( n140 ) ;
assign n142 =  ( slice_stream_full ) == ( 1'd1 )  ;
assign n143 =  ( n142 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n144 =  ( n39 ) ? ( LB2D_shift_7 ) : ( LB2D_shift_7 ) ;
assign n145 =  ( n34 ) ? ( LB2D_shift_7 ) : ( n144 ) ;
assign n146 =  ( n29 ) ? ( n143 ) : ( n145 ) ;
assign n147 =  ( n20 ) ? ( LB2D_shift_7 ) : ( n146 ) ;
assign n148 =  ( n11 ) ? ( LB2D_shift_7 ) : ( n147 ) ;
assign n149 =  ( n6 ) ? ( LB2D_shift_7 ) : ( n148 ) ;
assign n150 =  ( LB2D_shift_x ) == ( 9'd488 )  ;
assign n151 =  ( n21 ) & ( n150 )  ;
assign n152 =  ( n24 ) | ( n25 )  ;
assign n153 =  ( n151 ) & ( n152 )  ;
assign n154 =  ( LB2D_shift_x ) + ( 9'd1 )  ;
assign n155 =  ( n39 ) ? ( LB2D_shift_x ) : ( LB2D_shift_x ) ;
assign n156 =  ( n34 ) ? ( LB2D_shift_x ) : ( n155 ) ;
assign n157 =  ( n29 ) ? ( n154 ) : ( n156 ) ;
assign n158 =  ( n153 ) ? ( 9'd0 ) : ( n157 ) ;
assign n159 =  ( n20 ) ? ( LB2D_shift_x ) : ( n158 ) ;
assign n160 =  ( n11 ) ? ( LB2D_shift_x ) : ( n159 ) ;
assign n161 =  ( n6 ) ? ( LB2D_shift_x ) : ( n160 ) ;
assign n162 =  ( LB2D_shift_y ) < ( 10'd640 )  ;
assign n163 =  ( LB2D_shift_x ) < ( 9'd488 )  ;
assign n164 =  ( LB2D_shift_y ) + ( 10'd1 )  ;
assign n165 =  ( n163 ) ? ( LB2D_shift_y ) : ( n164 ) ;
assign n166 =  ( n162 ) ? ( n165 ) : ( 10'd640 ) ;
assign n167 =  ( n39 ) ? ( LB2D_shift_y ) : ( LB2D_shift_y ) ;
assign n168 =  ( n34 ) ? ( LB2D_shift_y ) : ( n167 ) ;
assign n169 =  ( n29 ) ? ( n166 ) : ( n168 ) ;
assign n170 =  ( n20 ) ? ( LB2D_shift_y ) : ( n169 ) ;
assign n171 =  ( n11 ) ? ( LB2D_shift_y ) : ( n170 ) ;
assign n172 =  ( n6 ) ? ( LB2D_shift_y ) : ( n171 ) ;
assign n173 =  ( stencil_stream_full ) == ( 1'd1 )  ;
assign n174 =  ( n173 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_0 ) ;
assign n175 = gb_fun(n174) ;
assign n176 =  ( n39 ) ? ( arg_0_TDATA ) : ( arg_0_TDATA ) ;
assign n177 =  ( n34 ) ? ( arg_0_TDATA ) : ( n176 ) ;
assign n178 =  ( n29 ) ? ( arg_0_TDATA ) : ( n177 ) ;
assign n179 =  ( n20 ) ? ( n175 ) : ( n178 ) ;
assign n180 =  ( n11 ) ? ( arg_0_TDATA ) : ( n179 ) ;
assign n181 =  ( n6 ) ? ( arg_0_TDATA ) : ( n180 ) ;
assign n182 =  ( gb_pp_it_8 ) == ( 1'd1 )  ;
assign n183 =  ( n182 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n184 =  ( n39 ) ? ( arg_0_TVALID ) : ( arg_0_TVALID ) ;
assign n185 =  ( n34 ) ? ( arg_0_TVALID ) : ( n184 ) ;
assign n186 =  ( n29 ) ? ( arg_0_TVALID ) : ( n185 ) ;
assign n187 =  ( n20 ) ? ( n183 ) : ( n186 ) ;
assign n188 =  ( n11 ) ? ( 1'd0 ) : ( n187 ) ;
assign n189 =  ( n6 ) ? ( arg_0_TVALID ) : ( n188 ) ;
assign n190 =  ( n39 ) ? ( 1'd1 ) : ( arg_1_TREADY ) ;
assign n191 =  ( n38 ) ? ( 1'd1 ) : ( n190 ) ;
assign n192 =  ( n34 ) ? ( arg_1_TREADY ) : ( n191 ) ;
assign n193 =  ( n29 ) ? ( arg_1_TREADY ) : ( n192 ) ;
assign n194 =  ( n20 ) ? ( arg_1_TREADY ) : ( n193 ) ;
assign n195 =  ( n11 ) ? ( arg_1_TREADY ) : ( n194 ) ;
assign n196 =  ( n6 ) ? ( 1'd1 ) : ( n195 ) ;
assign n197 =  ( gb_p_cnt ) == ( 19'd307200 )  ;
assign n198 =  ( n197 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n199 =  ( n39 ) ? ( gb_exit_it_1 ) : ( gb_exit_it_1 ) ;
assign n200 =  ( n34 ) ? ( gb_exit_it_1 ) : ( n199 ) ;
assign n201 =  ( n29 ) ? ( gb_exit_it_1 ) : ( n200 ) ;
assign n202 =  ( n20 ) ? ( n198 ) : ( n201 ) ;
assign n203 =  ( n11 ) ? ( gb_exit_it_1 ) : ( n202 ) ;
assign n204 =  ( n6 ) ? ( gb_exit_it_1 ) : ( n203 ) ;
assign n205 =  ( n39 ) ? ( gb_exit_it_2 ) : ( gb_exit_it_2 ) ;
assign n206 =  ( n34 ) ? ( gb_exit_it_2 ) : ( n205 ) ;
assign n207 =  ( n29 ) ? ( gb_exit_it_2 ) : ( n206 ) ;
assign n208 =  ( n20 ) ? ( gb_exit_it_1 ) : ( n207 ) ;
assign n209 =  ( n11 ) ? ( gb_exit_it_2 ) : ( n208 ) ;
assign n210 =  ( n6 ) ? ( gb_exit_it_2 ) : ( n209 ) ;
assign n211 =  ( n39 ) ? ( gb_exit_it_3 ) : ( gb_exit_it_3 ) ;
assign n212 =  ( n34 ) ? ( gb_exit_it_3 ) : ( n211 ) ;
assign n213 =  ( n29 ) ? ( gb_exit_it_3 ) : ( n212 ) ;
assign n214 =  ( n20 ) ? ( gb_exit_it_2 ) : ( n213 ) ;
assign n215 =  ( n11 ) ? ( gb_exit_it_3 ) : ( n214 ) ;
assign n216 =  ( n6 ) ? ( gb_exit_it_3 ) : ( n215 ) ;
assign n217 =  ( n39 ) ? ( gb_exit_it_4 ) : ( gb_exit_it_4 ) ;
assign n218 =  ( n34 ) ? ( gb_exit_it_4 ) : ( n217 ) ;
assign n219 =  ( n29 ) ? ( gb_exit_it_4 ) : ( n218 ) ;
assign n220 =  ( n20 ) ? ( gb_exit_it_3 ) : ( n219 ) ;
assign n221 =  ( n11 ) ? ( gb_exit_it_4 ) : ( n220 ) ;
assign n222 =  ( n6 ) ? ( gb_exit_it_4 ) : ( n221 ) ;
assign n223 =  ( n39 ) ? ( gb_exit_it_5 ) : ( gb_exit_it_5 ) ;
assign n224 =  ( n34 ) ? ( gb_exit_it_5 ) : ( n223 ) ;
assign n225 =  ( n29 ) ? ( gb_exit_it_5 ) : ( n224 ) ;
assign n226 =  ( n20 ) ? ( gb_exit_it_4 ) : ( n225 ) ;
assign n227 =  ( n11 ) ? ( gb_exit_it_5 ) : ( n226 ) ;
assign n228 =  ( n6 ) ? ( gb_exit_it_5 ) : ( n227 ) ;
assign n229 =  ( n39 ) ? ( gb_exit_it_6 ) : ( gb_exit_it_6 ) ;
assign n230 =  ( n34 ) ? ( gb_exit_it_6 ) : ( n229 ) ;
assign n231 =  ( n29 ) ? ( gb_exit_it_6 ) : ( n230 ) ;
assign n232 =  ( n20 ) ? ( gb_exit_it_5 ) : ( n231 ) ;
assign n233 =  ( n11 ) ? ( gb_exit_it_6 ) : ( n232 ) ;
assign n234 =  ( n6 ) ? ( gb_exit_it_6 ) : ( n233 ) ;
assign n235 =  ( n39 ) ? ( gb_exit_it_7 ) : ( gb_exit_it_7 ) ;
assign n236 =  ( n34 ) ? ( gb_exit_it_7 ) : ( n235 ) ;
assign n237 =  ( n29 ) ? ( gb_exit_it_7 ) : ( n236 ) ;
assign n238 =  ( n20 ) ? ( gb_exit_it_6 ) : ( n237 ) ;
assign n239 =  ( n11 ) ? ( gb_exit_it_7 ) : ( n238 ) ;
assign n240 =  ( n6 ) ? ( gb_exit_it_7 ) : ( n239 ) ;
assign n241 =  ( n39 ) ? ( gb_exit_it_8 ) : ( gb_exit_it_8 ) ;
assign n242 =  ( n34 ) ? ( gb_exit_it_8 ) : ( n241 ) ;
assign n243 =  ( n29 ) ? ( gb_exit_it_8 ) : ( n242 ) ;
assign n244 =  ( n20 ) ? ( gb_exit_it_7 ) : ( n243 ) ;
assign n245 =  ( n11 ) ? ( gb_exit_it_8 ) : ( n244 ) ;
assign n246 =  ( n6 ) ? ( gb_exit_it_8 ) : ( n245 ) ;
assign n247 =  ( gb_p_cnt ) < ( 19'd307200 )  ;
assign n248 =  ( gb_p_cnt ) + ( 19'd1 )  ;
assign n249 =  ( n247 ) ? ( n248 ) : ( 19'd307200 ) ;
assign n250 =  ( n39 ) ? ( gb_p_cnt ) : ( gb_p_cnt ) ;
assign n251 =  ( n34 ) ? ( gb_p_cnt ) : ( n250 ) ;
assign n252 =  ( n29 ) ? ( gb_p_cnt ) : ( n251 ) ;
assign n253 =  ( n20 ) ? ( n249 ) : ( n252 ) ;
assign n254 =  ( n11 ) ? ( gb_p_cnt ) : ( n253 ) ;
assign n255 =  ( n6 ) ? ( gb_p_cnt ) : ( n254 ) ;
assign n256 =  ( n39 ) ? ( gb_pp_it_1 ) : ( gb_pp_it_1 ) ;
assign n257 =  ( n34 ) ? ( gb_pp_it_1 ) : ( n256 ) ;
assign n258 =  ( n29 ) ? ( gb_pp_it_1 ) : ( n257 ) ;
assign n259 =  ( n20 ) ? ( 1'd1 ) : ( n258 ) ;
assign n260 =  ( n11 ) ? ( gb_pp_it_1 ) : ( n259 ) ;
assign n261 =  ( n6 ) ? ( gb_pp_it_1 ) : ( n260 ) ;
assign n262 =  ( n39 ) ? ( gb_pp_it_2 ) : ( gb_pp_it_2 ) ;
assign n263 =  ( n34 ) ? ( gb_pp_it_2 ) : ( n262 ) ;
assign n264 =  ( n29 ) ? ( gb_pp_it_2 ) : ( n263 ) ;
assign n265 =  ( n20 ) ? ( gb_pp_it_1 ) : ( n264 ) ;
assign n266 =  ( n11 ) ? ( gb_pp_it_2 ) : ( n265 ) ;
assign n267 =  ( n6 ) ? ( gb_pp_it_2 ) : ( n266 ) ;
assign n268 =  ( n39 ) ? ( gb_pp_it_3 ) : ( gb_pp_it_3 ) ;
assign n269 =  ( n34 ) ? ( gb_pp_it_3 ) : ( n268 ) ;
assign n270 =  ( n29 ) ? ( gb_pp_it_3 ) : ( n269 ) ;
assign n271 =  ( n20 ) ? ( gb_pp_it_2 ) : ( n270 ) ;
assign n272 =  ( n11 ) ? ( gb_pp_it_3 ) : ( n271 ) ;
assign n273 =  ( n6 ) ? ( gb_pp_it_3 ) : ( n272 ) ;
assign n274 =  ( n39 ) ? ( gb_pp_it_4 ) : ( gb_pp_it_4 ) ;
assign n275 =  ( n34 ) ? ( gb_pp_it_4 ) : ( n274 ) ;
assign n276 =  ( n29 ) ? ( gb_pp_it_4 ) : ( n275 ) ;
assign n277 =  ( n20 ) ? ( gb_pp_it_3 ) : ( n276 ) ;
assign n278 =  ( n11 ) ? ( gb_pp_it_4 ) : ( n277 ) ;
assign n279 =  ( n6 ) ? ( gb_pp_it_4 ) : ( n278 ) ;
assign n280 =  ( n39 ) ? ( gb_pp_it_5 ) : ( gb_pp_it_5 ) ;
assign n281 =  ( n34 ) ? ( gb_pp_it_5 ) : ( n280 ) ;
assign n282 =  ( n29 ) ? ( gb_pp_it_5 ) : ( n281 ) ;
assign n283 =  ( n20 ) ? ( gb_pp_it_4 ) : ( n282 ) ;
assign n284 =  ( n11 ) ? ( gb_pp_it_5 ) : ( n283 ) ;
assign n285 =  ( n6 ) ? ( gb_pp_it_5 ) : ( n284 ) ;
assign n286 =  ( n39 ) ? ( gb_pp_it_6 ) : ( gb_pp_it_6 ) ;
assign n287 =  ( n34 ) ? ( gb_pp_it_6 ) : ( n286 ) ;
assign n288 =  ( n29 ) ? ( gb_pp_it_6 ) : ( n287 ) ;
assign n289 =  ( n20 ) ? ( gb_pp_it_5 ) : ( n288 ) ;
assign n290 =  ( n11 ) ? ( gb_pp_it_6 ) : ( n289 ) ;
assign n291 =  ( n6 ) ? ( gb_pp_it_6 ) : ( n290 ) ;
assign n292 =  ( n39 ) ? ( gb_pp_it_7 ) : ( gb_pp_it_7 ) ;
assign n293 =  ( n34 ) ? ( gb_pp_it_7 ) : ( n292 ) ;
assign n294 =  ( n29 ) ? ( gb_pp_it_7 ) : ( n293 ) ;
assign n295 =  ( n20 ) ? ( gb_pp_it_6 ) : ( n294 ) ;
assign n296 =  ( n11 ) ? ( gb_pp_it_7 ) : ( n295 ) ;
assign n297 =  ( n6 ) ? ( gb_pp_it_7 ) : ( n296 ) ;
assign n298 =  ( n39 ) ? ( gb_pp_it_8 ) : ( gb_pp_it_8 ) ;
assign n299 =  ( n34 ) ? ( gb_pp_it_8 ) : ( n298 ) ;
assign n300 =  ( n29 ) ? ( gb_pp_it_8 ) : ( n299 ) ;
assign n301 =  ( n20 ) ? ( gb_pp_it_7 ) : ( n300 ) ;
assign n302 =  ( n11 ) ? ( gb_pp_it_8 ) : ( n301 ) ;
assign n303 =  ( n6 ) ? ( gb_pp_it_8 ) : ( n302 ) ;
assign n304 =  ( n39 ) ? ( gb_pp_it_9 ) : ( gb_pp_it_9 ) ;
assign n305 =  ( n34 ) ? ( gb_pp_it_9 ) : ( n304 ) ;
assign n306 =  ( n29 ) ? ( gb_pp_it_9 ) : ( n305 ) ;
assign n307 =  ( n20 ) ? ( gb_pp_it_8 ) : ( n306 ) ;
assign n308 =  ( n11 ) ? ( gb_pp_it_9 ) : ( n307 ) ;
assign n309 =  ( n6 ) ? ( gb_pp_it_9 ) : ( n308 ) ;
assign n310 =  ( n39 ) ? ( LB1D_uIn ) : ( in_stream_buff_0 ) ;
assign n311 =  ( n34 ) ? ( in_stream_buff_0 ) : ( n310 ) ;
assign n312 =  ( n29 ) ? ( in_stream_buff_0 ) : ( n311 ) ;
assign n313 =  ( n20 ) ? ( in_stream_buff_0 ) : ( n312 ) ;
assign n314 =  ( n11 ) ? ( in_stream_buff_0 ) : ( n313 ) ;
assign n315 =  ( n6 ) ? ( LB1D_uIn ) : ( n314 ) ;
assign n316 =  ( n39 ) ? ( in_stream_buff_0 ) : ( in_stream_buff_1 ) ;
assign n317 =  ( n34 ) ? ( in_stream_buff_1 ) : ( n316 ) ;
assign n318 =  ( n29 ) ? ( in_stream_buff_1 ) : ( n317 ) ;
assign n319 =  ( n20 ) ? ( in_stream_buff_1 ) : ( n318 ) ;
assign n320 =  ( n11 ) ? ( in_stream_buff_1 ) : ( n319 ) ;
assign n321 =  ( n6 ) ? ( in_stream_buff_0 ) : ( n320 ) ;
assign n322 =  ( in_stream_full ) == ( 1'd1 )  ;
assign n323 =  ( n322 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n324 =  ( n39 ) ? ( 1'd0 ) : ( in_stream_empty ) ;
assign n325 =  ( n34 ) ? ( n323 ) : ( n324 ) ;
assign n326 =  ( n29 ) ? ( in_stream_empty ) : ( n325 ) ;
assign n327 =  ( n20 ) ? ( in_stream_empty ) : ( n326 ) ;
assign n328 =  ( n11 ) ? ( in_stream_empty ) : ( n327 ) ;
assign n329 =  ( n6 ) ? ( 1'd0 ) : ( n328 ) ;
assign n330 =  ( in_stream_empty ) == ( 1'd1 )  ;
assign n331 =  ( n330 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n332 =  ( n39 ) ? ( n331 ) : ( in_stream_full ) ;
assign n333 =  ( n34 ) ? ( 1'd0 ) : ( n332 ) ;
assign n334 =  ( n29 ) ? ( in_stream_full ) : ( n333 ) ;
assign n335 =  ( n20 ) ? ( in_stream_full ) : ( n334 ) ;
assign n336 =  ( n11 ) ? ( in_stream_full ) : ( n335 ) ;
assign n337 =  ( n6 ) ? ( n331 ) : ( n336 ) ;
assign n338 =  ( n322 ) ? ( in_stream_buff_1 ) : ( in_stream_buff_0 ) ;
assign n339 =  ( LB2D_proc_w ) == ( 64'd0 )  ;
assign n340 =  ( LB2D_proc_x ) - ( 9'd1 )  ;
assign n341 =  (  LB2D_proc_7 [ n340 ] )  ;
assign n342 =  ( LB2D_proc_w ) == ( 64'd1 )  ;
assign n343 =  (  LB2D_proc_0 [ n340 ] )  ;
assign n344 =  ( LB2D_proc_w ) == ( 64'd2 )  ;
assign n345 =  (  LB2D_proc_1 [ n340 ] )  ;
assign n346 =  ( LB2D_proc_w ) == ( 64'd3 )  ;
assign n347 =  (  LB2D_proc_2 [ n340 ] )  ;
assign n348 =  ( LB2D_proc_w ) == ( 64'd4 )  ;
assign n349 =  (  LB2D_proc_3 [ n340 ] )  ;
assign n350 =  ( LB2D_proc_w ) == ( 64'd5 )  ;
assign n351 =  (  LB2D_proc_4 [ n340 ] )  ;
assign n352 =  ( LB2D_proc_w ) == ( 64'd6 )  ;
assign n353 =  (  LB2D_proc_5 [ n340 ] )  ;
assign n354 =  (  LB2D_proc_6 [ n340 ] )  ;
assign n355 =  ( n352 ) ? ( n353 ) : ( n354 ) ;
assign n356 =  ( n350 ) ? ( n351 ) : ( n355 ) ;
assign n357 =  ( n348 ) ? ( n349 ) : ( n356 ) ;
assign n358 =  ( n346 ) ? ( n347 ) : ( n357 ) ;
assign n359 =  ( n344 ) ? ( n345 ) : ( n358 ) ;
assign n360 =  ( n342 ) ? ( n343 ) : ( n359 ) ;
assign n361 =  ( n339 ) ? ( n341 ) : ( n360 ) ;
assign n362 =  ( n352 ) ? ( n351 ) : ( n353 ) ;
assign n363 =  ( n350 ) ? ( n349 ) : ( n362 ) ;
assign n364 =  ( n348 ) ? ( n347 ) : ( n363 ) ;
assign n365 =  ( n346 ) ? ( n345 ) : ( n364 ) ;
assign n366 =  ( n344 ) ? ( n343 ) : ( n365 ) ;
assign n367 =  ( n342 ) ? ( n341 ) : ( n366 ) ;
assign n368 =  ( n339 ) ? ( n354 ) : ( n367 ) ;
assign n369 =  ( n352 ) ? ( n349 ) : ( n351 ) ;
assign n370 =  ( n350 ) ? ( n347 ) : ( n369 ) ;
assign n371 =  ( n348 ) ? ( n345 ) : ( n370 ) ;
assign n372 =  ( n346 ) ? ( n343 ) : ( n371 ) ;
assign n373 =  ( n344 ) ? ( n341 ) : ( n372 ) ;
assign n374 =  ( n342 ) ? ( n354 ) : ( n373 ) ;
assign n375 =  ( n339 ) ? ( n353 ) : ( n374 ) ;
assign n376 =  ( n352 ) ? ( n347 ) : ( n349 ) ;
assign n377 =  ( n350 ) ? ( n345 ) : ( n376 ) ;
assign n378 =  ( n348 ) ? ( n343 ) : ( n377 ) ;
assign n379 =  ( n346 ) ? ( n341 ) : ( n378 ) ;
assign n380 =  ( n344 ) ? ( n354 ) : ( n379 ) ;
assign n381 =  ( n342 ) ? ( n353 ) : ( n380 ) ;
assign n382 =  ( n339 ) ? ( n351 ) : ( n381 ) ;
assign n383 =  ( n352 ) ? ( n345 ) : ( n347 ) ;
assign n384 =  ( n350 ) ? ( n343 ) : ( n383 ) ;
assign n385 =  ( n348 ) ? ( n341 ) : ( n384 ) ;
assign n386 =  ( n346 ) ? ( n354 ) : ( n385 ) ;
assign n387 =  ( n344 ) ? ( n353 ) : ( n386 ) ;
assign n388 =  ( n342 ) ? ( n351 ) : ( n387 ) ;
assign n389 =  ( n339 ) ? ( n349 ) : ( n388 ) ;
assign n390 =  ( n352 ) ? ( n343 ) : ( n345 ) ;
assign n391 =  ( n350 ) ? ( n341 ) : ( n390 ) ;
assign n392 =  ( n348 ) ? ( n354 ) : ( n391 ) ;
assign n393 =  ( n346 ) ? ( n353 ) : ( n392 ) ;
assign n394 =  ( n344 ) ? ( n351 ) : ( n393 ) ;
assign n395 =  ( n342 ) ? ( n349 ) : ( n394 ) ;
assign n396 =  ( n339 ) ? ( n347 ) : ( n395 ) ;
assign n397 =  ( n352 ) ? ( n341 ) : ( n343 ) ;
assign n398 =  ( n350 ) ? ( n354 ) : ( n397 ) ;
assign n399 =  ( n348 ) ? ( n353 ) : ( n398 ) ;
assign n400 =  ( n346 ) ? ( n351 ) : ( n399 ) ;
assign n401 =  ( n344 ) ? ( n349 ) : ( n400 ) ;
assign n402 =  ( n342 ) ? ( n347 ) : ( n401 ) ;
assign n403 =  ( n339 ) ? ( n345 ) : ( n402 ) ;
assign n404 =  ( n352 ) ? ( n354 ) : ( n341 ) ;
assign n405 =  ( n350 ) ? ( n353 ) : ( n404 ) ;
assign n406 =  ( n348 ) ? ( n351 ) : ( n405 ) ;
assign n407 =  ( n346 ) ? ( n349 ) : ( n406 ) ;
assign n408 =  ( n344 ) ? ( n347 ) : ( n407 ) ;
assign n409 =  ( n342 ) ? ( n345 ) : ( n408 ) ;
assign n410 =  ( n339 ) ? ( n343 ) : ( n409 ) ;
assign n411 =  { ( n403 ) , ( n410 ) }  ;
assign n412 =  { ( n396 ) , ( n411 ) }  ;
assign n413 =  { ( n389 ) , ( n412 ) }  ;
assign n414 =  { ( n382 ) , ( n413 ) }  ;
assign n415 =  { ( n375 ) , ( n414 ) }  ;
assign n416 =  { ( n368 ) , ( n415 ) }  ;
assign n417 =  { ( n361 ) , ( n416 ) }  ;
assign n418 =  { ( n338 ) , ( n417 ) }  ;
assign n419 =  ( n32 ) ? ( slice_stream_buff_0 ) : ( n418 ) ;
assign n420 =  ( n39 ) ? ( slice_stream_buff_0 ) : ( slice_stream_buff_0 ) ;
assign n421 =  ( n34 ) ? ( n419 ) : ( n420 ) ;
assign n422 =  ( n29 ) ? ( slice_stream_buff_0 ) : ( n421 ) ;
assign n423 =  ( n20 ) ? ( slice_stream_buff_0 ) : ( n422 ) ;
assign n424 =  ( n11 ) ? ( slice_stream_buff_0 ) : ( n423 ) ;
assign n425 =  ( n6 ) ? ( slice_stream_buff_0 ) : ( n424 ) ;
assign n426 =  ( n32 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n427 =  ( n39 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_1 ) ;
assign n428 =  ( n34 ) ? ( n426 ) : ( n427 ) ;
assign n429 =  ( n29 ) ? ( slice_stream_buff_1 ) : ( n428 ) ;
assign n430 =  ( n20 ) ? ( slice_stream_buff_1 ) : ( n429 ) ;
assign n431 =  ( n11 ) ? ( slice_stream_buff_1 ) : ( n430 ) ;
assign n432 =  ( n6 ) ? ( slice_stream_buff_1 ) : ( n431 ) ;
assign n433 =  ( n142 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n434 =  ( n32 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n435 =  ( n39 ) ? ( slice_stream_empty ) : ( slice_stream_empty ) ;
assign n436 =  ( n34 ) ? ( n434 ) : ( n435 ) ;
assign n437 =  ( n29 ) ? ( n433 ) : ( n436 ) ;
assign n438 =  ( n20 ) ? ( slice_stream_empty ) : ( n437 ) ;
assign n439 =  ( n11 ) ? ( slice_stream_empty ) : ( n438 ) ;
assign n440 =  ( n6 ) ? ( slice_stream_empty ) : ( n439 ) ;
assign n441 =  ( slice_stream_empty ) == ( 1'd1 )  ;
assign n442 =  ( n441 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n443 =  ( n32 ) ? ( 1'd0 ) : ( n442 ) ;
assign n444 =  ( n39 ) ? ( slice_stream_full ) : ( slice_stream_full ) ;
assign n445 =  ( n34 ) ? ( n443 ) : ( n444 ) ;
assign n446 =  ( n29 ) ? ( 1'd0 ) : ( n445 ) ;
assign n447 =  ( n20 ) ? ( slice_stream_full ) : ( n446 ) ;
assign n448 =  ( n11 ) ? ( slice_stream_full ) : ( n447 ) ;
assign n449 =  ( n6 ) ? ( slice_stream_full ) : ( n448 ) ;
assign n450 =  ( LB2D_shift_x ) >= ( 9'd8 )  ;
assign n451 =  ( LB2D_shift_x ) == ( 9'd0 )  ;
assign n452 =  ( n450 ) | ( n451 )  ;
assign n453 = n143[71:64] ;
assign n454 = LB2D_shift_7[71:64] ;
assign n455 = LB2D_shift_6[71:64] ;
assign n456 = LB2D_shift_5[71:64] ;
assign n457 = LB2D_shift_4[71:64] ;
assign n458 = LB2D_shift_3[71:64] ;
assign n459 = LB2D_shift_2[71:64] ;
assign n460 = LB2D_shift_1[71:64] ;
assign n461 = LB2D_shift_0[71:64] ;
assign n462 =  { ( n460 ) , ( n461 ) }  ;
assign n463 =  { ( n459 ) , ( n462 ) }  ;
assign n464 =  { ( n458 ) , ( n463 ) }  ;
assign n465 =  { ( n457 ) , ( n464 ) }  ;
assign n466 =  { ( n456 ) , ( n465 ) }  ;
assign n467 =  { ( n455 ) , ( n466 ) }  ;
assign n468 =  { ( n454 ) , ( n467 ) }  ;
assign n469 =  { ( n453 ) , ( n468 ) }  ;
assign n470 = n143[63:56] ;
assign n471 = LB2D_shift_7[63:56] ;
assign n472 = LB2D_shift_6[63:56] ;
assign n473 = LB2D_shift_5[63:56] ;
assign n474 = LB2D_shift_4[63:56] ;
assign n475 = LB2D_shift_3[63:56] ;
assign n476 = LB2D_shift_2[63:56] ;
assign n477 = LB2D_shift_1[63:56] ;
assign n478 = LB2D_shift_0[63:56] ;
assign n479 =  { ( n477 ) , ( n478 ) }  ;
assign n480 =  { ( n476 ) , ( n479 ) }  ;
assign n481 =  { ( n475 ) , ( n480 ) }  ;
assign n482 =  { ( n474 ) , ( n481 ) }  ;
assign n483 =  { ( n473 ) , ( n482 ) }  ;
assign n484 =  { ( n472 ) , ( n483 ) }  ;
assign n485 =  { ( n471 ) , ( n484 ) }  ;
assign n486 =  { ( n470 ) , ( n485 ) }  ;
assign n487 = n143[55:48] ;
assign n488 = LB2D_shift_7[55:48] ;
assign n489 = LB2D_shift_6[55:48] ;
assign n490 = LB2D_shift_5[55:48] ;
assign n491 = LB2D_shift_4[55:48] ;
assign n492 = LB2D_shift_3[55:48] ;
assign n493 = LB2D_shift_2[55:48] ;
assign n494 = LB2D_shift_1[55:48] ;
assign n495 = LB2D_shift_0[55:48] ;
assign n496 =  { ( n494 ) , ( n495 ) }  ;
assign n497 =  { ( n493 ) , ( n496 ) }  ;
assign n498 =  { ( n492 ) , ( n497 ) }  ;
assign n499 =  { ( n491 ) , ( n498 ) }  ;
assign n500 =  { ( n490 ) , ( n499 ) }  ;
assign n501 =  { ( n489 ) , ( n500 ) }  ;
assign n502 =  { ( n488 ) , ( n501 ) }  ;
assign n503 =  { ( n487 ) , ( n502 ) }  ;
assign n504 = n143[47:40] ;
assign n505 = LB2D_shift_7[47:40] ;
assign n506 = LB2D_shift_6[47:40] ;
assign n507 = LB2D_shift_5[47:40] ;
assign n508 = LB2D_shift_4[47:40] ;
assign n509 = LB2D_shift_3[47:40] ;
assign n510 = LB2D_shift_2[47:40] ;
assign n511 = LB2D_shift_1[47:40] ;
assign n512 = LB2D_shift_0[47:40] ;
assign n513 =  { ( n511 ) , ( n512 ) }  ;
assign n514 =  { ( n510 ) , ( n513 ) }  ;
assign n515 =  { ( n509 ) , ( n514 ) }  ;
assign n516 =  { ( n508 ) , ( n515 ) }  ;
assign n517 =  { ( n507 ) , ( n516 ) }  ;
assign n518 =  { ( n506 ) , ( n517 ) }  ;
assign n519 =  { ( n505 ) , ( n518 ) }  ;
assign n520 =  { ( n504 ) , ( n519 ) }  ;
assign n521 = n143[39:32] ;
assign n522 = LB2D_shift_7[39:32] ;
assign n523 = LB2D_shift_6[39:32] ;
assign n524 = LB2D_shift_5[39:32] ;
assign n525 = LB2D_shift_4[39:32] ;
assign n526 = LB2D_shift_3[39:32] ;
assign n527 = LB2D_shift_2[39:32] ;
assign n528 = LB2D_shift_1[39:32] ;
assign n529 = LB2D_shift_0[39:32] ;
assign n530 =  { ( n528 ) , ( n529 ) }  ;
assign n531 =  { ( n527 ) , ( n530 ) }  ;
assign n532 =  { ( n526 ) , ( n531 ) }  ;
assign n533 =  { ( n525 ) , ( n532 ) }  ;
assign n534 =  { ( n524 ) , ( n533 ) }  ;
assign n535 =  { ( n523 ) , ( n534 ) }  ;
assign n536 =  { ( n522 ) , ( n535 ) }  ;
assign n537 =  { ( n521 ) , ( n536 ) }  ;
assign n538 = n143[31:24] ;
assign n539 = LB2D_shift_7[31:24] ;
assign n540 = LB2D_shift_6[31:24] ;
assign n541 = LB2D_shift_5[31:24] ;
assign n542 = LB2D_shift_4[31:24] ;
assign n543 = LB2D_shift_3[31:24] ;
assign n544 = LB2D_shift_2[31:24] ;
assign n545 = LB2D_shift_1[31:24] ;
assign n546 = LB2D_shift_0[31:24] ;
assign n547 =  { ( n545 ) , ( n546 ) }  ;
assign n548 =  { ( n544 ) , ( n547 ) }  ;
assign n549 =  { ( n543 ) , ( n548 ) }  ;
assign n550 =  { ( n542 ) , ( n549 ) }  ;
assign n551 =  { ( n541 ) , ( n550 ) }  ;
assign n552 =  { ( n540 ) , ( n551 ) }  ;
assign n553 =  { ( n539 ) , ( n552 ) }  ;
assign n554 =  { ( n538 ) , ( n553 ) }  ;
assign n555 = n143[23:16] ;
assign n556 = LB2D_shift_7[23:16] ;
assign n557 = LB2D_shift_6[23:16] ;
assign n558 = LB2D_shift_5[23:16] ;
assign n559 = LB2D_shift_4[23:16] ;
assign n560 = LB2D_shift_3[23:16] ;
assign n561 = LB2D_shift_2[23:16] ;
assign n562 = LB2D_shift_1[23:16] ;
assign n563 = LB2D_shift_0[23:16] ;
assign n564 =  { ( n562 ) , ( n563 ) }  ;
assign n565 =  { ( n561 ) , ( n564 ) }  ;
assign n566 =  { ( n560 ) , ( n565 ) }  ;
assign n567 =  { ( n559 ) , ( n566 ) }  ;
assign n568 =  { ( n558 ) , ( n567 ) }  ;
assign n569 =  { ( n557 ) , ( n568 ) }  ;
assign n570 =  { ( n556 ) , ( n569 ) }  ;
assign n571 =  { ( n555 ) , ( n570 ) }  ;
assign n572 = n143[15:8] ;
assign n573 = LB2D_shift_7[15:8] ;
assign n574 = LB2D_shift_6[15:8] ;
assign n575 = LB2D_shift_5[15:8] ;
assign n576 = LB2D_shift_4[15:8] ;
assign n577 = LB2D_shift_3[15:8] ;
assign n578 = LB2D_shift_2[15:8] ;
assign n579 = LB2D_shift_1[15:8] ;
assign n580 = LB2D_shift_0[15:8] ;
assign n581 =  { ( n579 ) , ( n580 ) }  ;
assign n582 =  { ( n578 ) , ( n581 ) }  ;
assign n583 =  { ( n577 ) , ( n582 ) }  ;
assign n584 =  { ( n576 ) , ( n583 ) }  ;
assign n585 =  { ( n575 ) , ( n584 ) }  ;
assign n586 =  { ( n574 ) , ( n585 ) }  ;
assign n587 =  { ( n573 ) , ( n586 ) }  ;
assign n588 =  { ( n572 ) , ( n587 ) }  ;
assign n589 = n143[7:0] ;
assign n590 = LB2D_shift_7[7:0] ;
assign n591 = LB2D_shift_6[7:0] ;
assign n592 = LB2D_shift_5[7:0] ;
assign n593 = LB2D_shift_4[7:0] ;
assign n594 = LB2D_shift_3[7:0] ;
assign n595 = LB2D_shift_2[7:0] ;
assign n596 = LB2D_shift_1[7:0] ;
assign n597 = LB2D_shift_0[7:0] ;
assign n598 =  { ( n596 ) , ( n597 ) }  ;
assign n599 =  { ( n595 ) , ( n598 ) }  ;
assign n600 =  { ( n594 ) , ( n599 ) }  ;
assign n601 =  { ( n593 ) , ( n600 ) }  ;
assign n602 =  { ( n592 ) , ( n601 ) }  ;
assign n603 =  { ( n591 ) , ( n602 ) }  ;
assign n604 =  { ( n590 ) , ( n603 ) }  ;
assign n605 =  { ( n589 ) , ( n604 ) }  ;
assign n606 =  { ( n588 ) , ( n605 ) }  ;
assign n607 =  { ( n571 ) , ( n606 ) }  ;
assign n608 =  { ( n554 ) , ( n607 ) }  ;
assign n609 =  { ( n537 ) , ( n608 ) }  ;
assign n610 =  { ( n520 ) , ( n609 ) }  ;
assign n611 =  { ( n503 ) , ( n610 ) }  ;
assign n612 =  { ( n486 ) , ( n611 ) }  ;
assign n613 =  { ( n469 ) , ( n612 ) }  ;
assign n614 =  ( n452 ) ? ( n613 ) : ( stencil_stream_buff_0 ) ;
assign n615 =  ( n39 ) ? ( stencil_stream_buff_0 ) : ( stencil_stream_buff_0 ) ;
assign n616 =  ( n34 ) ? ( stencil_stream_buff_0 ) : ( n615 ) ;
assign n617 =  ( n29 ) ? ( n614 ) : ( n616 ) ;
assign n618 =  ( n20 ) ? ( stencil_stream_buff_0 ) : ( n617 ) ;
assign n619 =  ( n11 ) ? ( stencil_stream_buff_0 ) : ( n618 ) ;
assign n620 =  ( n6 ) ? ( stencil_stream_buff_0 ) : ( n619 ) ;
assign n621 =  ( n39 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_1 ) ;
assign n622 =  ( n34 ) ? ( stencil_stream_buff_1 ) : ( n621 ) ;
assign n623 =  ( n29 ) ? ( stencil_stream_buff_0 ) : ( n622 ) ;
assign n624 =  ( n20 ) ? ( stencil_stream_buff_1 ) : ( n623 ) ;
assign n625 =  ( n11 ) ? ( stencil_stream_buff_1 ) : ( n624 ) ;
assign n626 =  ( n6 ) ? ( stencil_stream_buff_1 ) : ( n625 ) ;
assign n627 =  ( n173 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n628 = ~ ( n452 ) ;
assign n629 =  ( n628 ) ? ( stencil_stream_empty ) : ( 1'd0 ) ;
assign n630 =  ( n39 ) ? ( stencil_stream_empty ) : ( stencil_stream_empty ) ;
assign n631 =  ( n34 ) ? ( stencil_stream_empty ) : ( n630 ) ;
assign n632 =  ( n29 ) ? ( n629 ) : ( n631 ) ;
assign n633 =  ( n20 ) ? ( n627 ) : ( n632 ) ;
assign n634 =  ( n11 ) ? ( stencil_stream_empty ) : ( n633 ) ;
assign n635 =  ( n6 ) ? ( stencil_stream_empty ) : ( n634 ) ;
assign n636 =  ( n16 ) ? ( 1'd0 ) : ( 1'd0 ) ;
assign n637 =  ( stencil_stream_empty ) == ( 1'd1 )  ;
assign n638 =  ( n637 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n639 =  ( n628 ) ? ( stencil_stream_full ) : ( n638 ) ;
assign n640 =  ( n39 ) ? ( stencil_stream_full ) : ( stencil_stream_full ) ;
assign n641 =  ( n34 ) ? ( stencil_stream_full ) : ( n640 ) ;
assign n642 =  ( n29 ) ? ( n639 ) : ( n641 ) ;
assign n643 =  ( n20 ) ? ( n636 ) : ( n642 ) ;
assign n644 =  ( n11 ) ? ( stencil_stream_full ) : ( n643 ) ;
assign n645 =  ( n6 ) ? ( stencil_stream_full ) : ( n644 ) ;
assign n646 = ~ ( n6 ) ;
assign n647 = ~ ( n11 ) ;
assign n648 =  ( n646 ) & ( n647 )  ;
assign n649 = ~ ( n20 ) ;
assign n650 =  ( n648 ) & ( n649 )  ;
assign n651 = ~ ( n29 ) ;
assign n652 =  ( n650 ) & ( n651 )  ;
assign n653 = ~ ( n34 ) ;
assign n654 =  ( n652 ) & ( n653 )  ;
assign n655 = ~ ( n39 ) ;
assign n656 =  ( n654 ) & ( n655 )  ;
assign n657 =  ( n654 ) & ( n39 )  ;
assign n658 =  ( n652 ) & ( n34 )  ;
assign n659 = ~ ( n339 ) ;
assign n660 =  ( n658 ) & ( n659 )  ;
assign n661 =  ( n658 ) & ( n339 )  ;
assign n662 =  ( n650 ) & ( n29 )  ;
assign n663 =  ( n648 ) & ( n20 )  ;
assign n664 =  ( n646 ) & ( n11 )  ;
assign LB2D_proc_0_addr0 = n661 ? (n340) : (0);
assign LB2D_proc_0_data0 = n661 ? (n338) : (LB2D_proc_0[0]);
assign n665 = ~ ( n342 ) ;
assign n666 =  ( n658 ) & ( n665 )  ;
assign n667 =  ( n658 ) & ( n342 )  ;
assign LB2D_proc_1_addr0 = n667 ? (n340) : (0);
assign LB2D_proc_1_data0 = n667 ? (n338) : (LB2D_proc_1[0]);
assign n668 = ~ ( n344 ) ;
assign n669 =  ( n658 ) & ( n668 )  ;
assign n670 =  ( n658 ) & ( n344 )  ;
assign LB2D_proc_2_addr0 = n670 ? (n340) : (0);
assign LB2D_proc_2_data0 = n670 ? (n338) : (LB2D_proc_2[0]);
assign n671 = ~ ( n346 ) ;
assign n672 =  ( n658 ) & ( n671 )  ;
assign n673 =  ( n658 ) & ( n346 )  ;
assign LB2D_proc_3_addr0 = n673 ? (n340) : (0);
assign LB2D_proc_3_data0 = n673 ? (n338) : (LB2D_proc_3[0]);
assign n674 = ~ ( n348 ) ;
assign n675 =  ( n658 ) & ( n674 )  ;
assign n676 =  ( n658 ) & ( n348 )  ;
assign LB2D_proc_4_addr0 = n676 ? (n340) : (0);
assign LB2D_proc_4_data0 = n676 ? (n338) : (LB2D_proc_4[0]);
assign n677 = ~ ( n350 ) ;
assign n678 =  ( n658 ) & ( n677 )  ;
assign n679 =  ( n658 ) & ( n350 )  ;
assign LB2D_proc_5_addr0 = n679 ? (n340) : (0);
assign LB2D_proc_5_data0 = n679 ? (n338) : (LB2D_proc_5[0]);
assign n680 = ~ ( n352 ) ;
assign n681 =  ( n658 ) & ( n680 )  ;
assign n682 =  ( n658 ) & ( n352 )  ;
assign LB2D_proc_6_addr0 = n682 ? (n340) : (0);
assign LB2D_proc_6_data0 = n682 ? (n338) : (LB2D_proc_6[0]);
assign n683 = ~ ( n72 ) ;
assign n684 =  ( n658 ) & ( n683 )  ;
assign n685 =  ( n658 ) & ( n72 )  ;
assign LB2D_proc_7_addr0 = n685 ? (n340) : (0);
assign LB2D_proc_7_data0 = n685 ? (n338) : (LB2D_proc_7[0]);
/*
function [7:0] gb_fun ;
input [647:0] arg0;
    begin
//TODO: Add the specific function HERE.    end
endfunction
*/

always @(posedge clk) begin
   if(rst) begin
       LB1D_buff <= LB1D_buff;
       LB1D_in <= LB1D_in;
       LB1D_it_1 <= LB1D_it_1;
       LB1D_p_cnt <= LB1D_p_cnt;
       LB1D_uIn <= LB1D_uIn;
       LB2D_proc_w <= LB2D_proc_w;
       LB2D_proc_x <= LB2D_proc_x;
       LB2D_proc_y <= LB2D_proc_y;
       LB2D_shift_0 <= LB2D_shift_0;
       LB2D_shift_1 <= LB2D_shift_1;
       LB2D_shift_2 <= LB2D_shift_2;
       LB2D_shift_3 <= LB2D_shift_3;
       LB2D_shift_4 <= LB2D_shift_4;
       LB2D_shift_5 <= LB2D_shift_5;
       LB2D_shift_6 <= LB2D_shift_6;
       LB2D_shift_7 <= LB2D_shift_7;
       LB2D_shift_x <= LB2D_shift_x;
       LB2D_shift_y <= LB2D_shift_y;
       arg_0_TDATA <= arg_0_TDATA;
       arg_0_TVALID <= arg_0_TVALID;
       arg_1_TREADY <= arg_1_TREADY;
       gb_exit_it_1 <= gb_exit_it_1;
       gb_exit_it_2 <= gb_exit_it_2;
       gb_exit_it_3 <= gb_exit_it_3;
       gb_exit_it_4 <= gb_exit_it_4;
       gb_exit_it_5 <= gb_exit_it_5;
       gb_exit_it_6 <= gb_exit_it_6;
       gb_exit_it_7 <= gb_exit_it_7;
       gb_exit_it_8 <= gb_exit_it_8;
       gb_p_cnt <= gb_p_cnt;
       gb_pp_it_1 <= gb_pp_it_1;
       gb_pp_it_2 <= gb_pp_it_2;
       gb_pp_it_3 <= gb_pp_it_3;
       gb_pp_it_4 <= gb_pp_it_4;
       gb_pp_it_5 <= gb_pp_it_5;
       gb_pp_it_6 <= gb_pp_it_6;
       gb_pp_it_7 <= gb_pp_it_7;
       gb_pp_it_8 <= gb_pp_it_8;
       gb_pp_it_9 <= gb_pp_it_9;
       in_stream_buff_0 <= in_stream_buff_0;
       in_stream_buff_1 <= in_stream_buff_1;
       in_stream_empty <= in_stream_empty;
       in_stream_full <= in_stream_full;
       slice_stream_buff_0 <= slice_stream_buff_0;
       slice_stream_buff_1 <= slice_stream_buff_1;
       slice_stream_empty <= slice_stream_empty;
       slice_stream_full <= slice_stream_full;
       stencil_stream_buff_0 <= stencil_stream_buff_0;
       stencil_stream_buff_1 <= stencil_stream_buff_1;
       stencil_stream_empty <= stencil_stream_empty;
       stencil_stream_full <= stencil_stream_full;
   end
   else if(step) begin
       LB1D_buff <= n46;
       LB1D_in <= n53;
       LB1D_it_1 <= n56;
       LB1D_p_cnt <= n64;
       LB1D_uIn <= n70;
       LB2D_proc_w <= n81;
       LB2D_proc_x <= n89;
       LB2D_proc_y <= n99;
       LB2D_shift_0 <= n105;
       LB2D_shift_1 <= n111;
       LB2D_shift_2 <= n117;
       LB2D_shift_3 <= n123;
       LB2D_shift_4 <= n129;
       LB2D_shift_5 <= n135;
       LB2D_shift_6 <= n141;
       LB2D_shift_7 <= n149;
       LB2D_shift_x <= n161;
       LB2D_shift_y <= n172;
       arg_0_TDATA <= n181;
       arg_0_TVALID <= n189;
       arg_1_TREADY <= n196;
       gb_exit_it_1 <= n204;
       gb_exit_it_2 <= n210;
       gb_exit_it_3 <= n216;
       gb_exit_it_4 <= n222;
       gb_exit_it_5 <= n228;
       gb_exit_it_6 <= n234;
       gb_exit_it_7 <= n240;
       gb_exit_it_8 <= n246;
       gb_p_cnt <= n255;
       gb_pp_it_1 <= n261;
       gb_pp_it_2 <= n267;
       gb_pp_it_3 <= n273;
       gb_pp_it_4 <= n279;
       gb_pp_it_5 <= n285;
       gb_pp_it_6 <= n291;
       gb_pp_it_7 <= n297;
       gb_pp_it_8 <= n303;
       gb_pp_it_9 <= n309;
       in_stream_buff_0 <= n315;
       in_stream_buff_1 <= n321;
       in_stream_empty <= n329;
       in_stream_full <= n337;
       slice_stream_buff_0 <= n425;
       slice_stream_buff_1 <= n432;
       slice_stream_empty <= n440;
       slice_stream_full <= n449;
       stencil_stream_buff_0 <= n620;
       stencil_stream_buff_1 <= n626;
       stencil_stream_empty <= n635;
       stencil_stream_full <= n645;
       LB2D_proc_0 [ LB2D_proc_0_addr0 ] <= LB2D_proc_0_data0;
       LB2D_proc_1 [ LB2D_proc_1_addr0 ] <= LB2D_proc_1_data0;
       LB2D_proc_2 [ LB2D_proc_2_addr0 ] <= LB2D_proc_2_data0;
       LB2D_proc_3 [ LB2D_proc_3_addr0 ] <= LB2D_proc_3_data0;
       LB2D_proc_4 [ LB2D_proc_4_addr0 ] <= LB2D_proc_4_data0;
       LB2D_proc_5 [ LB2D_proc_5_addr0 ] <= LB2D_proc_5_data0;
       LB2D_proc_6 [ LB2D_proc_6_addr0 ] <= LB2D_proc_6_data0;
       LB2D_proc_7 [ LB2D_proc_7_addr0 ] <= LB2D_proc_7_data0;
   end
end
endmodule
