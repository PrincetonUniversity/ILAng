module SPEC_B(
arg_0_TREADY,
arg_1_TDATA,
arg_1_TVALID,
LB1D_buff,
LB1D_in,
LB1D_it_1,
LB1D_p_cnt,
LB1D_uIn,
LB2D_proc_w,
LB2D_proc_x,
LB2D_proc_y,
LB2D_shift_0,
LB2D_shift_1,
LB2D_shift_2,
LB2D_shift_3,
LB2D_shift_4,
LB2D_shift_5,
LB2D_shift_6,
LB2D_shift_7,
LB2D_shift_x,
LB2D_shift_y,
arg_0_TDATA,
arg_0_TVALID,
arg_1_TREADY,
gb_exit_it_1,
gb_exit_it_2,
gb_exit_it_3,
gb_exit_it_4,
gb_exit_it_5,
gb_exit_it_6,
gb_exit_it_7,
gb_exit_it_8,
gb_p_cnt,
gb_pp_it_1,
gb_pp_it_2,
gb_pp_it_3,
gb_pp_it_4,
gb_pp_it_5,
gb_pp_it_6,
gb_pp_it_7,
gb_pp_it_8,
gb_pp_it_9,
in_stream_buff_0,
in_stream_buff_1,
in_stream_empty,
in_stream_full,
slice_stream_buff_0,
slice_stream_buff_1,
slice_stream_empty,
slice_stream_full,
stencil_stream_buff_0,
stencil_stream_buff_1,
stencil_stream_empty,
stencil_stream_full,
clk,rst,
step
);
input            arg_0_TREADY;
input      [7:0] arg_1_TDATA;
input            arg_1_TVALID;
input clk;
input rst;
input step;
output      [7:0] LB1D_buff;
output      [7:0] LB1D_in;
output            LB1D_it_1;
output     [18:0] LB1D_p_cnt;
output      [7:0] LB1D_uIn;
output     [63:0] LB2D_proc_w;
output      [8:0] LB2D_proc_x;
output      [9:0] LB2D_proc_y;
output     [71:0] LB2D_shift_0;
output     [71:0] LB2D_shift_1;
output     [71:0] LB2D_shift_2;
output     [71:0] LB2D_shift_3;
output     [71:0] LB2D_shift_4;
output     [71:0] LB2D_shift_5;
output     [71:0] LB2D_shift_6;
output     [71:0] LB2D_shift_7;
output      [8:0] LB2D_shift_x;
output      [9:0] LB2D_shift_y;
output      [7:0] arg_0_TDATA;
output            arg_0_TVALID;
output            arg_1_TREADY;
output            gb_exit_it_1;
output            gb_exit_it_2;
output            gb_exit_it_3;
output            gb_exit_it_4;
output            gb_exit_it_5;
output            gb_exit_it_6;
output            gb_exit_it_7;
output            gb_exit_it_8;
output     [18:0] gb_p_cnt;
output            gb_pp_it_1;
output            gb_pp_it_2;
output            gb_pp_it_3;
output            gb_pp_it_4;
output            gb_pp_it_5;
output            gb_pp_it_6;
output            gb_pp_it_7;
output            gb_pp_it_8;
output            gb_pp_it_9;
output      [7:0] in_stream_buff_0;
output      [7:0] in_stream_buff_1;
output            in_stream_empty;
output            in_stream_full;
output     [71:0] slice_stream_buff_0;
output     [71:0] slice_stream_buff_1;
output            slice_stream_empty;
output            slice_stream_full;
output    [647:0] stencil_stream_buff_0;
output    [647:0] stencil_stream_buff_1;
output            stencil_stream_empty;
output            stencil_stream_full;
reg      [7:0] LB1D_buff;
reg      [7:0] LB1D_in;
reg            LB1D_it_1;
reg     [18:0] LB1D_p_cnt;
reg      [7:0] LB1D_uIn;
reg     [63:0] LB2D_proc_w;
reg      [8:0] LB2D_proc_x;
reg      [9:0] LB2D_proc_y;
reg     [71:0] LB2D_shift_0;
reg     [71:0] LB2D_shift_1;
reg     [71:0] LB2D_shift_2;
reg     [71:0] LB2D_shift_3;
reg     [71:0] LB2D_shift_4;
reg     [71:0] LB2D_shift_5;
reg     [71:0] LB2D_shift_6;
reg     [71:0] LB2D_shift_7;
reg      [8:0] LB2D_shift_x;
reg      [9:0] LB2D_shift_y;
reg      [7:0] arg_0_TDATA;
reg            arg_0_TVALID;
reg            arg_1_TREADY;
reg            gb_exit_it_1;
reg            gb_exit_it_2;
reg            gb_exit_it_3;
reg            gb_exit_it_4;
reg            gb_exit_it_5;
reg            gb_exit_it_6;
reg            gb_exit_it_7;
reg            gb_exit_it_8;
reg     [18:0] gb_p_cnt;
reg            gb_pp_it_1;
reg            gb_pp_it_2;
reg            gb_pp_it_3;
reg            gb_pp_it_4;
reg            gb_pp_it_5;
reg            gb_pp_it_6;
reg            gb_pp_it_7;
reg            gb_pp_it_8;
reg            gb_pp_it_9;
reg      [7:0] in_stream_buff_0;
reg      [7:0] in_stream_buff_1;
reg            in_stream_empty;
reg            in_stream_full;
reg     [71:0] slice_stream_buff_0;
reg     [71:0] slice_stream_buff_1;
reg            slice_stream_empty;
reg            slice_stream_full;
reg    [647:0] stencil_stream_buff_0;
reg    [647:0] stencil_stream_buff_1;
reg            stencil_stream_empty;
reg            stencil_stream_full;
wire            arg_0_TREADY;
wire      [7:0] arg_1_TDATA;
wire            arg_1_TVALID;
wire            n0;
wire            n1;
wire            n2;
wire            n3;
wire            n4;
wire            n5;
wire            n6;
wire            n7;
wire            n8;
wire            n9;
wire            n10;
wire            n11;
wire            n12;
wire            n13;
wire            n14;
wire            n15;
wire            n16;
wire            n17;
wire            n18;
wire            n19;
wire            n20;
wire            n21;
wire            n22;
wire            n23;
wire            n24;
wire            n25;
wire            n26;
wire            n27;
wire            n28;
wire            n29;
wire            n30;
wire            n31;
wire            n32;
wire            n33;
wire            n34;
wire      [7:0] n35;
wire      [7:0] n36;
wire      [7:0] n37;
wire      [7:0] n38;
wire      [7:0] n39;
wire      [7:0] n40;
wire      [7:0] n41;
wire      [7:0] n42;
wire      [7:0] n43;
wire      [7:0] n44;
wire      [7:0] n45;
wire      [7:0] n46;
wire            n47;
wire            n48;
wire            n49;
wire            n50;
wire     [18:0] n51;
wire     [18:0] n52;
wire     [18:0] n53;
wire     [18:0] n54;
wire     [18:0] n55;
wire     [18:0] n56;
wire     [18:0] n57;
wire     [18:0] n58;
wire      [7:0] n59;
wire      [7:0] n60;
wire      [7:0] n61;
wire      [7:0] n62;
wire      [7:0] n63;
wire      [7:0] n64;
wire            n65;
wire            n66;
wire     [63:0] n67;
wire     [63:0] n68;
wire     [63:0] n69;
wire     [63:0] n70;
wire     [63:0] n71;
wire     [63:0] n72;
wire     [63:0] n73;
wire     [63:0] n74;
wire      [8:0] n75;
wire      [8:0] n76;
wire      [8:0] n77;
wire      [8:0] n78;
wire      [8:0] n79;
wire      [8:0] n80;
wire      [8:0] n81;
wire            n82;
wire      [9:0] n83;
wire      [9:0] n84;
wire      [9:0] n85;
wire      [9:0] n86;
wire      [9:0] n87;
wire      [9:0] n88;
wire      [9:0] n89;
wire      [9:0] n90;
wire     [71:0] n91;
wire     [71:0] n92;
wire     [71:0] n93;
wire     [71:0] n94;
wire     [71:0] n95;
wire     [71:0] n96;
wire     [71:0] n97;
wire     [71:0] n98;
wire     [71:0] n99;
wire     [71:0] n100;
wire     [71:0] n101;
wire     [71:0] n102;
wire     [71:0] n103;
wire     [71:0] n104;
wire     [71:0] n105;
wire     [71:0] n106;
wire     [71:0] n107;
wire     [71:0] n108;
wire     [71:0] n109;
wire     [71:0] n110;
wire     [71:0] n111;
wire     [71:0] n112;
wire     [71:0] n113;
wire     [71:0] n114;
wire     [71:0] n115;
wire     [71:0] n116;
wire     [71:0] n117;
wire     [71:0] n118;
wire     [71:0] n119;
wire     [71:0] n120;
wire     [71:0] n121;
wire     [71:0] n122;
wire     [71:0] n123;
wire     [71:0] n124;
wire     [71:0] n125;
wire            n126;
wire     [71:0] n127;
wire     [71:0] n128;
wire     [71:0] n129;
wire     [71:0] n130;
wire     [71:0] n131;
wire     [71:0] n132;
wire            n133;
wire            n134;
wire            n135;
wire            n136;
wire      [8:0] n137;
wire      [8:0] n138;
wire      [8:0] n139;
wire      [8:0] n140;
wire      [8:0] n141;
wire      [8:0] n142;
wire      [8:0] n143;
wire            n144;
wire            n145;
wire      [9:0] n146;
wire      [9:0] n147;
wire      [9:0] n148;
wire      [9:0] n149;
wire      [9:0] n150;
wire      [9:0] n151;
wire      [9:0] n152;
wire      [9:0] n153;
wire            n154;
wire    [647:0] n155;
wire      [7:0] n156;
wire      [7:0] n157;
wire      [7:0] n158;
wire      [7:0] n159;
wire      [7:0] n160;
wire      [7:0] n161;
wire            n162;
wire            n163;
wire            n164;
wire            n165;
wire            n166;
wire            n167;
wire            n168;
wire     [18:0] n169;
wire            n170;
wire            n171;
wire            n172;
wire            n173;
wire            n174;
wire            n175;
wire            n176;
wire            n177;
wire     [18:0] n178;
wire            n179;
wire            n180;
wire            n181;
wire            n182;
wire            n183;
wire            n184;
wire            n185;
wire            n186;
wire            n187;
wire            n188;
wire            n189;
wire            n190;
wire            n191;
wire            n192;
wire            n193;
wire            n194;
wire            n195;
wire            n196;
wire            n197;
wire            n198;
wire            n199;
wire            n200;
wire            n201;
wire            n202;
wire            n203;
wire            n204;
wire            n205;
wire            n206;
wire            n207;
wire            n208;
wire            n209;
wire            n210;
wire            n211;
wire            n212;
wire            n213;
wire            n214;
wire            n215;
wire            n216;
wire            n217;
wire            n218;
wire            n219;
wire            n220;
wire            n221;
wire     [18:0] n222;
wire     [18:0] n223;
wire     [18:0] n224;
wire     [18:0] n225;
wire     [18:0] n226;
wire     [18:0] n227;
wire            n228;
wire            n229;
wire            n230;
wire            n231;
wire            n232;
wire            n233;
wire            n234;
wire            n235;
wire            n236;
wire            n237;
wire            n238;
wire            n239;
wire            n240;
wire            n241;
wire            n242;
wire            n243;
wire            n244;
wire            n245;
wire            n246;
wire            n247;
wire            n248;
wire            n249;
wire            n250;
wire            n251;
wire            n252;
wire            n253;
wire            n254;
wire            n255;
wire            n256;
wire            n257;
wire            n258;
wire            n259;
wire            n260;
wire            n261;
wire            n262;
wire            n263;
wire            n264;
wire            n265;
wire            n266;
wire            n267;
wire            n268;
wire            n269;
wire            n270;
wire            n271;
wire            n272;
wire      [7:0] n273;
wire      [7:0] n274;
wire      [7:0] n275;
wire      [7:0] n276;
wire      [7:0] n277;
wire      [7:0] n278;
wire      [7:0] n279;
wire      [7:0] n280;
wire      [7:0] n281;
wire      [7:0] n282;
wire            n283;
wire            n284;
wire            n285;
wire            n286;
wire            n287;
wire            n288;
wire            n289;
wire            n290;
wire            n291;
wire            n292;
wire            n293;
wire            n294;
wire            n295;
wire            n296;
wire      [7:0] n297;
wire            n298;
wire      [8:0] n299;
wire      [7:0] n300;
wire            n301;
wire      [7:0] n302;
wire            n303;
wire      [7:0] n304;
wire            n305;
wire      [7:0] n306;
wire            n307;
wire      [7:0] n308;
wire            n309;
wire      [7:0] n310;
wire            n311;
wire      [7:0] n312;
wire      [7:0] n313;
wire      [7:0] n314;
wire      [7:0] n315;
wire      [7:0] n316;
wire      [7:0] n317;
wire      [7:0] n318;
wire      [7:0] n319;
wire      [7:0] n320;
wire      [7:0] n321;
wire      [7:0] n322;
wire      [7:0] n323;
wire      [7:0] n324;
wire      [7:0] n325;
wire      [7:0] n326;
wire      [7:0] n327;
wire      [7:0] n328;
wire      [7:0] n329;
wire      [7:0] n330;
wire      [7:0] n331;
wire      [7:0] n332;
wire      [7:0] n333;
wire      [7:0] n334;
wire      [7:0] n335;
wire      [7:0] n336;
wire      [7:0] n337;
wire      [7:0] n338;
wire      [7:0] n339;
wire      [7:0] n340;
wire      [7:0] n341;
wire      [7:0] n342;
wire      [7:0] n343;
wire      [7:0] n344;
wire      [7:0] n345;
wire      [7:0] n346;
wire      [7:0] n347;
wire      [7:0] n348;
wire      [7:0] n349;
wire      [7:0] n350;
wire      [7:0] n351;
wire      [7:0] n352;
wire      [7:0] n353;
wire      [7:0] n354;
wire      [7:0] n355;
wire      [7:0] n356;
wire      [7:0] n357;
wire      [7:0] n358;
wire      [7:0] n359;
wire      [7:0] n360;
wire      [7:0] n361;
wire      [7:0] n362;
wire      [7:0] n363;
wire      [7:0] n364;
wire      [7:0] n365;
wire      [7:0] n366;
wire      [7:0] n367;
wire      [7:0] n368;
wire      [7:0] n369;
wire     [15:0] n370;
wire     [23:0] n371;
wire     [31:0] n372;
wire     [39:0] n373;
wire     [47:0] n374;
wire     [55:0] n375;
wire     [63:0] n376;
wire     [71:0] n377;
wire     [71:0] n378;
wire     [71:0] n379;
wire     [71:0] n380;
wire     [71:0] n381;
wire     [71:0] n382;
wire     [71:0] n383;
wire     [71:0] n384;
wire     [71:0] n385;
wire     [71:0] n386;
wire     [71:0] n387;
wire     [71:0] n388;
wire     [71:0] n389;
wire            n390;
wire            n391;
wire            n392;
wire            n393;
wire            n394;
wire            n395;
wire            n396;
wire            n397;
wire            n398;
wire            n399;
wire            n400;
wire            n401;
wire            n402;
wire            n403;
wire            n404;
wire            n405;
wire            n406;
wire            n407;
wire      [7:0] n408;
wire      [7:0] n409;
wire      [7:0] n410;
wire      [7:0] n411;
wire      [7:0] n412;
wire      [7:0] n413;
wire      [7:0] n414;
wire      [7:0] n415;
wire      [7:0] n416;
wire     [15:0] n417;
wire     [23:0] n418;
wire     [31:0] n419;
wire     [39:0] n420;
wire     [47:0] n421;
wire     [55:0] n422;
wire     [63:0] n423;
wire     [71:0] n424;
wire      [7:0] n425;
wire      [7:0] n426;
wire      [7:0] n427;
wire      [7:0] n428;
wire      [7:0] n429;
wire      [7:0] n430;
wire      [7:0] n431;
wire      [7:0] n432;
wire      [7:0] n433;
wire     [15:0] n434;
wire     [23:0] n435;
wire     [31:0] n436;
wire     [39:0] n437;
wire     [47:0] n438;
wire     [55:0] n439;
wire     [63:0] n440;
wire     [71:0] n441;
wire      [7:0] n442;
wire      [7:0] n443;
wire      [7:0] n444;
wire      [7:0] n445;
wire      [7:0] n446;
wire      [7:0] n447;
wire      [7:0] n448;
wire      [7:0] n449;
wire      [7:0] n450;
wire     [15:0] n451;
wire     [23:0] n452;
wire     [31:0] n453;
wire     [39:0] n454;
wire     [47:0] n455;
wire     [55:0] n456;
wire     [63:0] n457;
wire     [71:0] n458;
wire      [7:0] n459;
wire      [7:0] n460;
wire      [7:0] n461;
wire      [7:0] n462;
wire      [7:0] n463;
wire      [7:0] n464;
wire      [7:0] n465;
wire      [7:0] n466;
wire      [7:0] n467;
wire     [15:0] n468;
wire     [23:0] n469;
wire     [31:0] n470;
wire     [39:0] n471;
wire     [47:0] n472;
wire     [55:0] n473;
wire     [63:0] n474;
wire     [71:0] n475;
wire      [7:0] n476;
wire      [7:0] n477;
wire      [7:0] n478;
wire      [7:0] n479;
wire      [7:0] n480;
wire      [7:0] n481;
wire      [7:0] n482;
wire      [7:0] n483;
wire      [7:0] n484;
wire     [15:0] n485;
wire     [23:0] n486;
wire     [31:0] n487;
wire     [39:0] n488;
wire     [47:0] n489;
wire     [55:0] n490;
wire     [63:0] n491;
wire     [71:0] n492;
wire      [7:0] n493;
wire      [7:0] n494;
wire      [7:0] n495;
wire      [7:0] n496;
wire      [7:0] n497;
wire      [7:0] n498;
wire      [7:0] n499;
wire      [7:0] n500;
wire      [7:0] n501;
wire     [15:0] n502;
wire     [23:0] n503;
wire     [31:0] n504;
wire     [39:0] n505;
wire     [47:0] n506;
wire     [55:0] n507;
wire     [63:0] n508;
wire     [71:0] n509;
wire      [7:0] n510;
wire      [7:0] n511;
wire      [7:0] n512;
wire      [7:0] n513;
wire      [7:0] n514;
wire      [7:0] n515;
wire      [7:0] n516;
wire      [7:0] n517;
wire      [7:0] n518;
wire     [15:0] n519;
wire     [23:0] n520;
wire     [31:0] n521;
wire     [39:0] n522;
wire     [47:0] n523;
wire     [55:0] n524;
wire     [63:0] n525;
wire     [71:0] n526;
wire      [7:0] n527;
wire      [7:0] n528;
wire      [7:0] n529;
wire      [7:0] n530;
wire      [7:0] n531;
wire      [7:0] n532;
wire      [7:0] n533;
wire      [7:0] n534;
wire      [7:0] n535;
wire     [15:0] n536;
wire     [23:0] n537;
wire     [31:0] n538;
wire     [39:0] n539;
wire     [47:0] n540;
wire     [55:0] n541;
wire     [63:0] n542;
wire     [71:0] n543;
wire      [7:0] n544;
wire      [7:0] n545;
wire      [7:0] n546;
wire      [7:0] n547;
wire      [7:0] n548;
wire      [7:0] n549;
wire      [7:0] n550;
wire      [7:0] n551;
wire      [7:0] n552;
wire     [15:0] n553;
wire     [23:0] n554;
wire     [31:0] n555;
wire     [39:0] n556;
wire     [47:0] n557;
wire     [55:0] n558;
wire     [63:0] n559;
wire     [71:0] n560;
wire    [143:0] n561;
wire    [215:0] n562;
wire    [287:0] n563;
wire    [359:0] n564;
wire    [431:0] n565;
wire    [503:0] n566;
wire    [575:0] n567;
wire    [647:0] n568;
wire    [647:0] n569;
wire    [647:0] n570;
wire    [647:0] n571;
wire    [647:0] n572;
wire    [647:0] n573;
wire    [647:0] n574;
wire    [647:0] n575;
wire    [647:0] n576;
wire    [647:0] n577;
wire    [647:0] n578;
wire    [647:0] n579;
wire            n580;
wire            n581;
wire            n582;
wire            n583;
wire            n584;
wire            n585;
wire            n586;
wire            n587;
wire            n588;
wire            n589;
wire            n590;
wire            n591;
wire            n592;
wire            n593;
wire            n594;
wire            n595;
wire            n596;
wire      [8:0] LB2D_proc_0_addr0;
wire      [7:0] LB2D_proc_0_data0;
wire            n597;
wire            n598;
wire            n599;
wire            n600;
wire            n601;
wire            n602;
wire            n603;
wire            n604;
wire            n605;
wire            n606;
wire            n607;
wire            n608;
wire            n609;
wire            n610;
wire            n611;
wire            n612;
wire      [8:0] LB2D_proc_1_addr0;
wire      [7:0] LB2D_proc_1_data0;
wire            n613;
wire            n614;
wire            n615;
wire      [8:0] LB2D_proc_2_addr0;
wire      [7:0] LB2D_proc_2_data0;
wire            n616;
wire            n617;
wire            n618;
wire      [8:0] LB2D_proc_3_addr0;
wire      [7:0] LB2D_proc_3_data0;
wire            n619;
wire            n620;
wire            n621;
wire      [8:0] LB2D_proc_4_addr0;
wire      [7:0] LB2D_proc_4_data0;
wire            n622;
wire            n623;
wire            n624;
wire      [8:0] LB2D_proc_5_addr0;
wire      [7:0] LB2D_proc_5_data0;
wire            n625;
wire            n626;
wire            n627;
wire      [8:0] LB2D_proc_6_addr0;
wire      [7:0] LB2D_proc_6_data0;
wire            n628;
wire            n629;
wire            n630;
wire      [8:0] LB2D_proc_7_addr0;
wire      [7:0] LB2D_proc_7_data0;
wire            n631;
wire            n632;
wire            n633;
reg      [7:0] LB2D_proc_0[487:0];
reg      [7:0] LB2D_proc_1[487:0];
reg      [7:0] LB2D_proc_2[487:0];
reg      [7:0] LB2D_proc_3[487:0];
reg      [7:0] LB2D_proc_4[487:0];
reg      [7:0] LB2D_proc_5[487:0];
reg      [7:0] LB2D_proc_6[487:0];
reg      [7:0] LB2D_proc_7[487:0];
wire clk;
wire rst;
wire step;
assign n0 =  ( arg_1_TREADY ) == ( 1'd1 )  ;
assign n1 =  ( arg_1_TVALID ) == ( 1'd1 )  ;
assign n2 =  ( n0 ) & ( n1 )  ;
assign n3 =  ( arg_0_TREADY ) == ( 1'd0 )  ;
assign n4 =  ( n2 ) & ( n3 )  ;
assign n5 =  ( arg_0_TVALID ) == ( 1'd0 )  ;
assign n6 =  ( gb_exit_it_1 ) == ( 1'd0 )  ;
assign n7 =  ( stencil_stream_empty ) == ( 1'd0 )  ;
assign n8 =  ( n6 ) & ( n7 )  ;
assign n9 =  ( gb_exit_it_1 ) == ( 1'd1 )  ;
assign n10 =  ( gb_exit_it_8 ) == ( 1'd0 )  ;
assign n11 =  ( n9 ) & ( n10 )  ;
assign n12 =  ( n8 ) | ( n11 )  ;
assign n13 =  ( n5 ) & ( n12 )  ;
assign n14 =  ( slice_stream_empty ) == ( 1'd0 )  ;
assign n15 =  ( LB2D_shift_x ) != ( 9'd488 )  ;
assign n16 =  ( n14 ) & ( n15 )  ;
assign n17 =  ( stencil_stream_full ) == ( 1'd0 )  ;
assign n18 =  ( LB2D_shift_x ) < ( 9'd8 )  ;
assign n19 =  ( LB2D_shift_x ) > ( 9'd0 )  ;
assign n20 =  ( n18 ) & ( n19 )  ;
assign n21 =  ( n17 ) | ( n20 )  ;
assign n22 =  ( n16 ) & ( n21 )  ;
assign n23 =  ( in_stream_empty ) == ( 1'd0 )  ;
assign n24 =  ( slice_stream_full ) == ( 1'd0 )  ;
assign n25 =  ( LB2D_proc_y ) < ( 10'd8 )  ;
assign n26 =  ( n24 ) | ( n25 )  ;
assign n27 =  ( n23 ) & ( n26 )  ;
assign n28 =  ( arg_1_TREADY ) == ( 1'd0 )  ;
assign n29 =  ( in_stream_full ) == ( 1'd0 )  ;
assign n30 =  ( n28 ) & ( n29 )  ;
assign n31 =  ( LB1D_it_1 ) == ( 1'd0 )  ;
assign n32 =  ( n30 ) & ( n31 )  ;
assign n33 =  ( LB1D_it_1 ) == ( 1'd1 )  ;
assign n34 =  ( n30 ) & ( n33 )  ;
assign n35 =  ( n34 ) ? ( LB1D_uIn ) : ( LB1D_buff ) ;
assign n36 =  ( n32 ) ? ( LB1D_uIn ) : ( n35 ) ;
assign n37 =  ( n27 ) ? ( LB1D_buff ) : ( n36 ) ;
assign n38 =  ( n22 ) ? ( LB1D_buff ) : ( n37 ) ;
assign n39 =  ( n13 ) ? ( LB1D_buff ) : ( n38 ) ;
assign n40 =  ( n4 ) ? ( LB1D_buff ) : ( n39 ) ;
assign n41 =  ( n34 ) ? ( LB1D_in ) : ( LB1D_in ) ;
assign n42 =  ( n32 ) ? ( LB1D_in ) : ( n41 ) ;
assign n43 =  ( n27 ) ? ( LB1D_in ) : ( n42 ) ;
assign n44 =  ( n22 ) ? ( LB1D_in ) : ( n43 ) ;
assign n45 =  ( n13 ) ? ( LB1D_in ) : ( n44 ) ;
assign n46 =  ( n4 ) ? ( arg_1_TDATA ) : ( n45 ) ;
assign n47 =  ( LB1D_p_cnt ) == ( 19'd316224 )  ;
assign n48 =  ( n47 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n49 =  ( n34 ) ? ( n48 ) : ( LB1D_it_1 ) ;
assign n50 =  ( n32 ) ? ( 1'd1 ) : ( n49 ) ;
assign n51 =  ( LB1D_p_cnt ) + ( 19'd1 )  ;
assign n52 =  ( n47 ) ? ( 19'd0 ) : ( n51 ) ;
assign n53 =  ( n34 ) ? ( n52 ) : ( LB1D_p_cnt ) ;
assign n54 =  ( n32 ) ? ( n51 ) : ( n53 ) ;
assign n55 =  ( n27 ) ? ( LB1D_p_cnt ) : ( n54 ) ;
assign n56 =  ( n22 ) ? ( LB1D_p_cnt ) : ( n55 ) ;
assign n57 =  ( n13 ) ? ( LB1D_p_cnt ) : ( n56 ) ;
assign n58 =  ( n4 ) ? ( LB1D_p_cnt ) : ( n57 ) ;
assign n59 =  ( n34 ) ? ( LB1D_in ) : ( LB1D_uIn ) ;
assign n60 =  ( n32 ) ? ( LB1D_in ) : ( n59 ) ;
assign n61 =  ( n27 ) ? ( LB1D_uIn ) : ( n60 ) ;
assign n62 =  ( n22 ) ? ( LB1D_uIn ) : ( n61 ) ;
assign n63 =  ( n13 ) ? ( LB1D_uIn ) : ( n62 ) ;
assign n64 =  ( n4 ) ? ( LB1D_uIn ) : ( n63 ) ;
assign n65 =  ( LB2D_proc_x ) == ( 9'd488 )  ;
assign n66 =  ( LB2D_proc_w ) == ( 64'd7 )  ;
assign n67 =  ( LB2D_proc_w ) + ( 64'd1 )  ;
assign n68 =  ( n66 ) ? ( 64'd0 ) : ( n67 ) ;
assign n69 =  ( n65 ) ? ( n68 ) : ( LB2D_proc_w ) ;
assign n70 =  ( n34 ) ? ( LB2D_proc_w ) : ( LB2D_proc_w ) ;
assign n71 =  ( n27 ) ? ( n69 ) : ( n70 ) ;
assign n72 =  ( n22 ) ? ( LB2D_proc_w ) : ( n71 ) ;
assign n73 =  ( n13 ) ? ( LB2D_proc_w ) : ( n72 ) ;
assign n74 =  ( n4 ) ? ( LB2D_proc_w ) : ( n73 ) ;
assign n75 =  ( LB2D_proc_x ) + ( 9'd1 )  ;
assign n76 =  ( n65 ) ? ( 9'd1 ) : ( n75 ) ;
assign n77 =  ( n34 ) ? ( LB2D_proc_x ) : ( LB2D_proc_x ) ;
assign n78 =  ( n27 ) ? ( n76 ) : ( n77 ) ;
assign n79 =  ( n22 ) ? ( LB2D_proc_x ) : ( n78 ) ;
assign n80 =  ( n13 ) ? ( LB2D_proc_x ) : ( n79 ) ;
assign n81 =  ( n4 ) ? ( LB2D_proc_x ) : ( n80 ) ;
assign n82 =  ( LB2D_proc_y ) == ( 10'd648 )  ;
assign n83 =  ( LB2D_proc_y ) + ( 10'd1 )  ;
assign n84 =  ( n82 ) ? ( 10'd0 ) : ( n83 ) ;
assign n85 =  ( n65 ) ? ( n84 ) : ( LB2D_proc_y ) ;
assign n86 =  ( n34 ) ? ( LB2D_proc_y ) : ( LB2D_proc_y ) ;
assign n87 =  ( n27 ) ? ( n85 ) : ( n86 ) ;
assign n88 =  ( n22 ) ? ( LB2D_proc_y ) : ( n87 ) ;
assign n89 =  ( n13 ) ? ( LB2D_proc_y ) : ( n88 ) ;
assign n90 =  ( n4 ) ? ( LB2D_proc_y ) : ( n89 ) ;
assign n91 =  ( n34 ) ? ( LB2D_shift_0 ) : ( LB2D_shift_0 ) ;
assign n92 =  ( n27 ) ? ( LB2D_shift_0 ) : ( n91 ) ;
assign n93 =  ( n22 ) ? ( LB2D_shift_1 ) : ( n92 ) ;
assign n94 =  ( n13 ) ? ( LB2D_shift_0 ) : ( n93 ) ;
assign n95 =  ( n4 ) ? ( LB2D_shift_0 ) : ( n94 ) ;
assign n96 =  ( n34 ) ? ( LB2D_shift_1 ) : ( LB2D_shift_1 ) ;
assign n97 =  ( n27 ) ? ( LB2D_shift_1 ) : ( n96 ) ;
assign n98 =  ( n22 ) ? ( LB2D_shift_2 ) : ( n97 ) ;
assign n99 =  ( n13 ) ? ( LB2D_shift_1 ) : ( n98 ) ;
assign n100 =  ( n4 ) ? ( LB2D_shift_1 ) : ( n99 ) ;
assign n101 =  ( n34 ) ? ( LB2D_shift_2 ) : ( LB2D_shift_2 ) ;
assign n102 =  ( n27 ) ? ( LB2D_shift_2 ) : ( n101 ) ;
assign n103 =  ( n22 ) ? ( LB2D_shift_3 ) : ( n102 ) ;
assign n104 =  ( n13 ) ? ( LB2D_shift_2 ) : ( n103 ) ;
assign n105 =  ( n4 ) ? ( LB2D_shift_2 ) : ( n104 ) ;
assign n106 =  ( n34 ) ? ( LB2D_shift_3 ) : ( LB2D_shift_3 ) ;
assign n107 =  ( n27 ) ? ( LB2D_shift_3 ) : ( n106 ) ;
assign n108 =  ( n22 ) ? ( LB2D_shift_4 ) : ( n107 ) ;
assign n109 =  ( n13 ) ? ( LB2D_shift_3 ) : ( n108 ) ;
assign n110 =  ( n4 ) ? ( LB2D_shift_3 ) : ( n109 ) ;
assign n111 =  ( n34 ) ? ( LB2D_shift_4 ) : ( LB2D_shift_4 ) ;
assign n112 =  ( n27 ) ? ( LB2D_shift_4 ) : ( n111 ) ;
assign n113 =  ( n22 ) ? ( LB2D_shift_5 ) : ( n112 ) ;
assign n114 =  ( n13 ) ? ( LB2D_shift_4 ) : ( n113 ) ;
assign n115 =  ( n4 ) ? ( LB2D_shift_4 ) : ( n114 ) ;
assign n116 =  ( n34 ) ? ( LB2D_shift_5 ) : ( LB2D_shift_5 ) ;
assign n117 =  ( n27 ) ? ( LB2D_shift_5 ) : ( n116 ) ;
assign n118 =  ( n22 ) ? ( LB2D_shift_6 ) : ( n117 ) ;
assign n119 =  ( n13 ) ? ( LB2D_shift_5 ) : ( n118 ) ;
assign n120 =  ( n4 ) ? ( LB2D_shift_5 ) : ( n119 ) ;
assign n121 =  ( n34 ) ? ( LB2D_shift_6 ) : ( LB2D_shift_6 ) ;
assign n122 =  ( n27 ) ? ( LB2D_shift_6 ) : ( n121 ) ;
assign n123 =  ( n22 ) ? ( LB2D_shift_7 ) : ( n122 ) ;
assign n124 =  ( n13 ) ? ( LB2D_shift_6 ) : ( n123 ) ;
assign n125 =  ( n4 ) ? ( LB2D_shift_6 ) : ( n124 ) ;
assign n126 =  ( slice_stream_full ) == ( 1'd1 )  ;
assign n127 =  ( n126 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n128 =  ( n34 ) ? ( LB2D_shift_7 ) : ( LB2D_shift_7 ) ;
assign n129 =  ( n27 ) ? ( LB2D_shift_7 ) : ( n128 ) ;
assign n130 =  ( n22 ) ? ( n127 ) : ( n129 ) ;
assign n131 =  ( n13 ) ? ( LB2D_shift_7 ) : ( n130 ) ;
assign n132 =  ( n4 ) ? ( LB2D_shift_7 ) : ( n131 ) ;
assign n133 =  ( LB2D_shift_x ) == ( 9'd488 )  ;
assign n134 =  ( n14 ) & ( n133 )  ;
assign n135 =  ( n17 ) | ( n18 )  ;
assign n136 =  ( n134 ) & ( n135 )  ;
assign n137 =  ( LB2D_shift_x ) + ( 9'd1 )  ;
assign n138 =  ( n34 ) ? ( LB2D_shift_x ) : ( LB2D_shift_x ) ;
assign n139 =  ( n27 ) ? ( LB2D_shift_x ) : ( n138 ) ;
assign n140 =  ( n22 ) ? ( n137 ) : ( n139 ) ;
assign n141 =  ( n136 ) ? ( 9'd0 ) : ( n140 ) ;
assign n142 =  ( n13 ) ? ( LB2D_shift_x ) : ( n141 ) ;
assign n143 =  ( n4 ) ? ( LB2D_shift_x ) : ( n142 ) ;
assign n144 =  ( LB2D_shift_y ) < ( 10'd640 )  ;
assign n145 =  ( LB2D_shift_x ) < ( 9'd488 )  ;
assign n146 =  ( LB2D_shift_y ) + ( 10'd1 )  ;
assign n147 =  ( n145 ) ? ( LB2D_shift_y ) : ( n146 ) ;
assign n148 =  ( n144 ) ? ( n147 ) : ( 10'd640 ) ;
assign n149 =  ( n34 ) ? ( LB2D_shift_y ) : ( LB2D_shift_y ) ;
assign n150 =  ( n27 ) ? ( LB2D_shift_y ) : ( n149 ) ;
assign n151 =  ( n22 ) ? ( n148 ) : ( n150 ) ;
assign n152 =  ( n13 ) ? ( LB2D_shift_y ) : ( n151 ) ;
assign n153 =  ( n4 ) ? ( LB2D_shift_y ) : ( n152 ) ;
assign n154 =  ( stencil_stream_full ) == ( 1'd1 )  ;
assign n155 =  ( n154 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_0 ) ;
//assign n156 = gb_fun(n155) ;
gb_fun gb_fun_U (
        .a (n155),
        .b (n156)
        );

assign n157 =  ( n34 ) ? ( arg_0_TDATA ) : ( arg_0_TDATA ) ;
assign n158 =  ( n27 ) ? ( arg_0_TDATA ) : ( n157 ) ;
assign n159 =  ( n22 ) ? ( arg_0_TDATA ) : ( n158 ) ;
assign n160 =  ( n13 ) ? ( n156 ) : ( n159 ) ;
assign n161 =  ( n4 ) ? ( arg_0_TDATA ) : ( n160 ) ;
assign n162 =  ( gb_pp_it_8 ) == ( 1'd1 )  ;
assign n163 =  ( n162 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n164 =  ( n34 ) ? ( arg_0_TVALID ) : ( arg_0_TVALID ) ;
assign n165 =  ( n27 ) ? ( arg_0_TVALID ) : ( n164 ) ;
assign n166 =  ( n22 ) ? ( arg_0_TVALID ) : ( n165 ) ;
assign n167 =  ( n13 ) ? ( n163 ) : ( n166 ) ;
assign n168 =  ( n4 ) ? ( arg_0_TVALID ) : ( n167 ) ;
assign n169 =  ( 19'd316224 ) - ( 19'd1 )  ;
assign n170 =  ( LB1D_p_cnt ) == ( n169 )  ;
assign n171 =  ( n170 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n172 =  ( n34 ) ? ( n171 ) : ( arg_1_TREADY ) ;
assign n173 =  ( n32 ) ? ( 1'd1 ) : ( n172 ) ;
assign n174 =  ( n27 ) ? ( arg_1_TREADY ) : ( n173 ) ;
assign n175 =  ( n22 ) ? ( arg_1_TREADY ) : ( n174 ) ;
assign n176 =  ( n13 ) ? ( arg_1_TREADY ) : ( n175 ) ;
assign n177 =  ( n4 ) ? ( 1'd0 ) : ( n176 ) ;
assign n178 =  ( gb_p_cnt ) + ( 19'd1 )  ;
assign n179 =  ( n178 ) == ( 19'd307200 )  ;
assign n180 =  ( n179 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n181 =  ( n34 ) ? ( gb_exit_it_1 ) : ( gb_exit_it_1 ) ;
assign n182 =  ( n27 ) ? ( gb_exit_it_1 ) : ( n181 ) ;
assign n183 =  ( n22 ) ? ( gb_exit_it_1 ) : ( n182 ) ;
assign n184 =  ( n13 ) ? ( n180 ) : ( n183 ) ;
assign n185 =  ( n4 ) ? ( gb_exit_it_1 ) : ( n184 ) ;
assign n186 =  ( n34 ) ? ( gb_exit_it_2 ) : ( gb_exit_it_2 ) ;
assign n187 =  ( n27 ) ? ( gb_exit_it_2 ) : ( n186 ) ;
assign n188 =  ( n22 ) ? ( gb_exit_it_2 ) : ( n187 ) ;
assign n189 =  ( n13 ) ? ( gb_exit_it_1 ) : ( n188 ) ;
assign n190 =  ( n4 ) ? ( gb_exit_it_2 ) : ( n189 ) ;
assign n191 =  ( n34 ) ? ( gb_exit_it_3 ) : ( gb_exit_it_3 ) ;
assign n192 =  ( n27 ) ? ( gb_exit_it_3 ) : ( n191 ) ;
assign n193 =  ( n22 ) ? ( gb_exit_it_3 ) : ( n192 ) ;
assign n194 =  ( n13 ) ? ( gb_exit_it_2 ) : ( n193 ) ;
assign n195 =  ( n4 ) ? ( gb_exit_it_3 ) : ( n194 ) ;
assign n196 =  ( n34 ) ? ( gb_exit_it_4 ) : ( gb_exit_it_4 ) ;
assign n197 =  ( n27 ) ? ( gb_exit_it_4 ) : ( n196 ) ;
assign n198 =  ( n22 ) ? ( gb_exit_it_4 ) : ( n197 ) ;
assign n199 =  ( n13 ) ? ( gb_exit_it_3 ) : ( n198 ) ;
assign n200 =  ( n4 ) ? ( gb_exit_it_4 ) : ( n199 ) ;
assign n201 =  ( n34 ) ? ( gb_exit_it_5 ) : ( gb_exit_it_5 ) ;
assign n202 =  ( n27 ) ? ( gb_exit_it_5 ) : ( n201 ) ;
assign n203 =  ( n22 ) ? ( gb_exit_it_5 ) : ( n202 ) ;
assign n204 =  ( n13 ) ? ( gb_exit_it_4 ) : ( n203 ) ;
assign n205 =  ( n4 ) ? ( gb_exit_it_5 ) : ( n204 ) ;
assign n206 =  ( n34 ) ? ( gb_exit_it_6 ) : ( gb_exit_it_6 ) ;
assign n207 =  ( n27 ) ? ( gb_exit_it_6 ) : ( n206 ) ;
assign n208 =  ( n22 ) ? ( gb_exit_it_6 ) : ( n207 ) ;
assign n209 =  ( n13 ) ? ( gb_exit_it_5 ) : ( n208 ) ;
assign n210 =  ( n4 ) ? ( gb_exit_it_6 ) : ( n209 ) ;
assign n211 =  ( n34 ) ? ( gb_exit_it_7 ) : ( gb_exit_it_7 ) ;
assign n212 =  ( n27 ) ? ( gb_exit_it_7 ) : ( n211 ) ;
assign n213 =  ( n22 ) ? ( gb_exit_it_7 ) : ( n212 ) ;
assign n214 =  ( n13 ) ? ( gb_exit_it_6 ) : ( n213 ) ;
assign n215 =  ( n4 ) ? ( gb_exit_it_7 ) : ( n214 ) ;
assign n216 =  ( n34 ) ? ( gb_exit_it_8 ) : ( gb_exit_it_8 ) ;
assign n217 =  ( n27 ) ? ( gb_exit_it_8 ) : ( n216 ) ;
assign n218 =  ( n22 ) ? ( gb_exit_it_8 ) : ( n217 ) ;
assign n219 =  ( n13 ) ? ( gb_exit_it_7 ) : ( n218 ) ;
assign n220 =  ( n4 ) ? ( gb_exit_it_8 ) : ( n219 ) ;
assign n221 =  ( gb_p_cnt ) < ( 19'd307200 )  ;
assign n222 =  ( n221 ) ? ( n178 ) : ( 19'd307200 ) ;
assign n223 =  ( n34 ) ? ( gb_p_cnt ) : ( gb_p_cnt ) ;
assign n224 =  ( n27 ) ? ( gb_p_cnt ) : ( n223 ) ;
assign n225 =  ( n22 ) ? ( gb_p_cnt ) : ( n224 ) ;
assign n226 =  ( n13 ) ? ( n222 ) : ( n225 ) ;
assign n227 =  ( n4 ) ? ( gb_p_cnt ) : ( n226 ) ;
assign n228 =  ( n34 ) ? ( gb_pp_it_1 ) : ( gb_pp_it_1 ) ;
assign n229 =  ( n27 ) ? ( gb_pp_it_1 ) : ( n228 ) ;
assign n230 =  ( n22 ) ? ( gb_pp_it_1 ) : ( n229 ) ;
assign n231 =  ( n13 ) ? ( 1'd1 ) : ( n230 ) ;
assign n232 =  ( n4 ) ? ( gb_pp_it_1 ) : ( n231 ) ;
assign n233 =  ( n34 ) ? ( gb_pp_it_2 ) : ( gb_pp_it_2 ) ;
assign n234 =  ( n27 ) ? ( gb_pp_it_2 ) : ( n233 ) ;
assign n235 =  ( n22 ) ? ( gb_pp_it_2 ) : ( n234 ) ;
assign n236 =  ( n13 ) ? ( gb_pp_it_1 ) : ( n235 ) ;
assign n237 =  ( n4 ) ? ( gb_pp_it_2 ) : ( n236 ) ;
assign n238 =  ( n34 ) ? ( gb_pp_it_3 ) : ( gb_pp_it_3 ) ;
assign n239 =  ( n27 ) ? ( gb_pp_it_3 ) : ( n238 ) ;
assign n240 =  ( n22 ) ? ( gb_pp_it_3 ) : ( n239 ) ;
assign n241 =  ( n13 ) ? ( gb_pp_it_2 ) : ( n240 ) ;
assign n242 =  ( n4 ) ? ( gb_pp_it_3 ) : ( n241 ) ;
assign n243 =  ( n34 ) ? ( gb_pp_it_4 ) : ( gb_pp_it_4 ) ;
assign n244 =  ( n27 ) ? ( gb_pp_it_4 ) : ( n243 ) ;
assign n245 =  ( n22 ) ? ( gb_pp_it_4 ) : ( n244 ) ;
assign n246 =  ( n13 ) ? ( gb_pp_it_3 ) : ( n245 ) ;
assign n247 =  ( n4 ) ? ( gb_pp_it_4 ) : ( n246 ) ;
assign n248 =  ( n34 ) ? ( gb_pp_it_5 ) : ( gb_pp_it_5 ) ;
assign n249 =  ( n27 ) ? ( gb_pp_it_5 ) : ( n248 ) ;
assign n250 =  ( n22 ) ? ( gb_pp_it_5 ) : ( n249 ) ;
assign n251 =  ( n13 ) ? ( gb_pp_it_4 ) : ( n250 ) ;
assign n252 =  ( n4 ) ? ( gb_pp_it_5 ) : ( n251 ) ;
assign n253 =  ( n34 ) ? ( gb_pp_it_6 ) : ( gb_pp_it_6 ) ;
assign n254 =  ( n27 ) ? ( gb_pp_it_6 ) : ( n253 ) ;
assign n255 =  ( n22 ) ? ( gb_pp_it_6 ) : ( n254 ) ;
assign n256 =  ( n13 ) ? ( gb_pp_it_5 ) : ( n255 ) ;
assign n257 =  ( n4 ) ? ( gb_pp_it_6 ) : ( n256 ) ;
assign n258 =  ( n34 ) ? ( gb_pp_it_7 ) : ( gb_pp_it_7 ) ;
assign n259 =  ( n27 ) ? ( gb_pp_it_7 ) : ( n258 ) ;
assign n260 =  ( n22 ) ? ( gb_pp_it_7 ) : ( n259 ) ;
assign n261 =  ( n13 ) ? ( gb_pp_it_6 ) : ( n260 ) ;
assign n262 =  ( n4 ) ? ( gb_pp_it_7 ) : ( n261 ) ;
assign n263 =  ( n34 ) ? ( gb_pp_it_8 ) : ( gb_pp_it_8 ) ;
assign n264 =  ( n27 ) ? ( gb_pp_it_8 ) : ( n263 ) ;
assign n265 =  ( n22 ) ? ( gb_pp_it_8 ) : ( n264 ) ;
assign n266 =  ( n13 ) ? ( gb_pp_it_7 ) : ( n265 ) ;
assign n267 =  ( n4 ) ? ( gb_pp_it_8 ) : ( n266 ) ;
assign n268 =  ( n34 ) ? ( gb_pp_it_9 ) : ( gb_pp_it_9 ) ;
assign n269 =  ( n27 ) ? ( gb_pp_it_9 ) : ( n268 ) ;
assign n270 =  ( n22 ) ? ( gb_pp_it_9 ) : ( n269 ) ;
assign n271 =  ( n13 ) ? ( gb_pp_it_8 ) : ( n270 ) ;
assign n272 =  ( n4 ) ? ( gb_pp_it_9 ) : ( n271 ) ;
assign n273 =  ( n34 ) ? ( LB1D_buff ) : ( in_stream_buff_0 ) ;
assign n274 =  ( n27 ) ? ( in_stream_buff_0 ) : ( n273 ) ;
assign n275 =  ( n22 ) ? ( in_stream_buff_0 ) : ( n274 ) ;
assign n276 =  ( n13 ) ? ( in_stream_buff_0 ) : ( n275 ) ;
assign n277 =  ( n4 ) ? ( in_stream_buff_0 ) : ( n276 ) ;
assign n278 =  ( n34 ) ? ( in_stream_buff_0 ) : ( in_stream_buff_1 ) ;
assign n279 =  ( n27 ) ? ( in_stream_buff_1 ) : ( n278 ) ;
assign n280 =  ( n22 ) ? ( in_stream_buff_1 ) : ( n279 ) ;
assign n281 =  ( n13 ) ? ( in_stream_buff_1 ) : ( n280 ) ;
assign n282 =  ( n4 ) ? ( in_stream_buff_1 ) : ( n281 ) ;
assign n283 =  ( in_stream_full ) == ( 1'd1 )  ;
assign n284 =  ( n283 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n285 =  ( n34 ) ? ( 1'd0 ) : ( in_stream_empty ) ;
assign n286 =  ( n27 ) ? ( n284 ) : ( n285 ) ;
assign n287 =  ( n22 ) ? ( in_stream_empty ) : ( n286 ) ;
assign n288 =  ( n13 ) ? ( in_stream_empty ) : ( n287 ) ;
assign n289 =  ( n4 ) ? ( in_stream_empty ) : ( n288 ) ;
assign n290 =  ( in_stream_empty ) == ( 1'd1 )  ;
assign n291 =  ( n290 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n292 =  ( n34 ) ? ( n291 ) : ( in_stream_full ) ;
assign n293 =  ( n27 ) ? ( 1'd0 ) : ( n292 ) ;
assign n294 =  ( n22 ) ? ( in_stream_full ) : ( n293 ) ;
assign n295 =  ( n13 ) ? ( in_stream_full ) : ( n294 ) ;
assign n296 =  ( n4 ) ? ( in_stream_full ) : ( n295 ) ;
assign n297 =  ( n283 ) ? ( in_stream_buff_1 ) : ( in_stream_buff_0 ) ;
assign n298 =  ( LB2D_proc_w ) == ( 64'd0 )  ;
assign n299 =  ( LB2D_proc_x ) - ( 9'd1 )  ;
assign n300 =  (  LB2D_proc_7 [ n299 ] )  ;
assign n301 =  ( LB2D_proc_w ) == ( 64'd1 )  ;
assign n302 =  (  LB2D_proc_0 [ n299 ] )  ;
assign n303 =  ( LB2D_proc_w ) == ( 64'd2 )  ;
assign n304 =  (  LB2D_proc_1 [ n299 ] )  ;
assign n305 =  ( LB2D_proc_w ) == ( 64'd3 )  ;
assign n306 =  (  LB2D_proc_2 [ n299 ] )  ;
assign n307 =  ( LB2D_proc_w ) == ( 64'd4 )  ;
assign n308 =  (  LB2D_proc_3 [ n299 ] )  ;
assign n309 =  ( LB2D_proc_w ) == ( 64'd5 )  ;
assign n310 =  (  LB2D_proc_4 [ n299 ] )  ;
assign n311 =  ( LB2D_proc_w ) == ( 64'd6 )  ;
assign n312 =  (  LB2D_proc_5 [ n299 ] )  ;
assign n313 =  (  LB2D_proc_6 [ n299 ] )  ;
assign n314 =  ( n311 ) ? ( n312 ) : ( n313 ) ;
assign n315 =  ( n309 ) ? ( n310 ) : ( n314 ) ;
assign n316 =  ( n307 ) ? ( n308 ) : ( n315 ) ;
assign n317 =  ( n305 ) ? ( n306 ) : ( n316 ) ;
assign n318 =  ( n303 ) ? ( n304 ) : ( n317 ) ;
assign n319 =  ( n301 ) ? ( n302 ) : ( n318 ) ;
assign n320 =  ( n298 ) ? ( n300 ) : ( n319 ) ;
assign n321 =  ( n311 ) ? ( n310 ) : ( n312 ) ;
assign n322 =  ( n309 ) ? ( n308 ) : ( n321 ) ;
assign n323 =  ( n307 ) ? ( n306 ) : ( n322 ) ;
assign n324 =  ( n305 ) ? ( n304 ) : ( n323 ) ;
assign n325 =  ( n303 ) ? ( n302 ) : ( n324 ) ;
assign n326 =  ( n301 ) ? ( n300 ) : ( n325 ) ;
assign n327 =  ( n298 ) ? ( n313 ) : ( n326 ) ;
assign n328 =  ( n311 ) ? ( n308 ) : ( n310 ) ;
assign n329 =  ( n309 ) ? ( n306 ) : ( n328 ) ;
assign n330 =  ( n307 ) ? ( n304 ) : ( n329 ) ;
assign n331 =  ( n305 ) ? ( n302 ) : ( n330 ) ;
assign n332 =  ( n303 ) ? ( n300 ) : ( n331 ) ;
assign n333 =  ( n301 ) ? ( n313 ) : ( n332 ) ;
assign n334 =  ( n298 ) ? ( n312 ) : ( n333 ) ;
assign n335 =  ( n311 ) ? ( n306 ) : ( n308 ) ;
assign n336 =  ( n309 ) ? ( n304 ) : ( n335 ) ;
assign n337 =  ( n307 ) ? ( n302 ) : ( n336 ) ;
assign n338 =  ( n305 ) ? ( n300 ) : ( n337 ) ;
assign n339 =  ( n303 ) ? ( n313 ) : ( n338 ) ;
assign n340 =  ( n301 ) ? ( n312 ) : ( n339 ) ;
assign n341 =  ( n298 ) ? ( n310 ) : ( n340 ) ;
assign n342 =  ( n311 ) ? ( n304 ) : ( n306 ) ;
assign n343 =  ( n309 ) ? ( n302 ) : ( n342 ) ;
assign n344 =  ( n307 ) ? ( n300 ) : ( n343 ) ;
assign n345 =  ( n305 ) ? ( n313 ) : ( n344 ) ;
assign n346 =  ( n303 ) ? ( n312 ) : ( n345 ) ;
assign n347 =  ( n301 ) ? ( n310 ) : ( n346 ) ;
assign n348 =  ( n298 ) ? ( n308 ) : ( n347 ) ;
assign n349 =  ( n311 ) ? ( n302 ) : ( n304 ) ;
assign n350 =  ( n309 ) ? ( n300 ) : ( n349 ) ;
assign n351 =  ( n307 ) ? ( n313 ) : ( n350 ) ;
assign n352 =  ( n305 ) ? ( n312 ) : ( n351 ) ;
assign n353 =  ( n303 ) ? ( n310 ) : ( n352 ) ;
assign n354 =  ( n301 ) ? ( n308 ) : ( n353 ) ;
assign n355 =  ( n298 ) ? ( n306 ) : ( n354 ) ;
assign n356 =  ( n311 ) ? ( n300 ) : ( n302 ) ;
assign n357 =  ( n309 ) ? ( n313 ) : ( n356 ) ;
assign n358 =  ( n307 ) ? ( n312 ) : ( n357 ) ;
assign n359 =  ( n305 ) ? ( n310 ) : ( n358 ) ;
assign n360 =  ( n303 ) ? ( n308 ) : ( n359 ) ;
assign n361 =  ( n301 ) ? ( n306 ) : ( n360 ) ;
assign n362 =  ( n298 ) ? ( n304 ) : ( n361 ) ;
assign n363 =  ( n311 ) ? ( n313 ) : ( n300 ) ;
assign n364 =  ( n309 ) ? ( n312 ) : ( n363 ) ;
assign n365 =  ( n307 ) ? ( n310 ) : ( n364 ) ;
assign n366 =  ( n305 ) ? ( n308 ) : ( n365 ) ;
assign n367 =  ( n303 ) ? ( n306 ) : ( n366 ) ;
assign n368 =  ( n301 ) ? ( n304 ) : ( n367 ) ;
assign n369 =  ( n298 ) ? ( n302 ) : ( n368 ) ;
assign n370 =  { ( n362 ) , ( n369 ) }  ;
assign n371 =  { ( n355 ) , ( n370 ) }  ;
assign n372 =  { ( n348 ) , ( n371 ) }  ;
assign n373 =  { ( n341 ) , ( n372 ) }  ;
assign n374 =  { ( n334 ) , ( n373 ) }  ;
assign n375 =  { ( n327 ) , ( n374 ) }  ;
assign n376 =  { ( n320 ) , ( n375 ) }  ;
assign n377 =  { ( n297 ) , ( n376 ) }  ;
assign n378 =  ( n25 ) ? ( slice_stream_buff_0 ) : ( n377 ) ;
assign n379 =  ( n34 ) ? ( slice_stream_buff_0 ) : ( slice_stream_buff_0 ) ;
assign n380 =  ( n27 ) ? ( n378 ) : ( n379 ) ;
assign n381 =  ( n22 ) ? ( slice_stream_buff_0 ) : ( n380 ) ;
assign n382 =  ( n13 ) ? ( slice_stream_buff_0 ) : ( n381 ) ;
assign n383 =  ( n4 ) ? ( slice_stream_buff_0 ) : ( n382 ) ;
assign n384 =  ( n25 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n385 =  ( n34 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_1 ) ;
assign n386 =  ( n27 ) ? ( n384 ) : ( n385 ) ;
assign n387 =  ( n22 ) ? ( slice_stream_buff_1 ) : ( n386 ) ;
assign n388 =  ( n13 ) ? ( slice_stream_buff_1 ) : ( n387 ) ;
assign n389 =  ( n4 ) ? ( slice_stream_buff_1 ) : ( n388 ) ;
assign n390 =  ( n126 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n391 =  ( n25 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n392 =  ( n34 ) ? ( slice_stream_empty ) : ( slice_stream_empty ) ;
assign n393 =  ( n27 ) ? ( n391 ) : ( n392 ) ;
assign n394 =  ( n22 ) ? ( n390 ) : ( n393 ) ;
assign n395 =  ( n13 ) ? ( slice_stream_empty ) : ( n394 ) ;
assign n396 =  ( n4 ) ? ( slice_stream_empty ) : ( n395 ) ;
assign n397 =  ( slice_stream_empty ) == ( 1'd1 )  ;
assign n398 =  ( n397 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n399 =  ( n25 ) ? ( 1'd0 ) : ( n398 ) ;
assign n400 =  ( n34 ) ? ( slice_stream_full ) : ( slice_stream_full ) ;
assign n401 =  ( n27 ) ? ( n399 ) : ( n400 ) ;
assign n402 =  ( n22 ) ? ( 1'd0 ) : ( n401 ) ;
assign n403 =  ( n13 ) ? ( slice_stream_full ) : ( n402 ) ;
assign n404 =  ( n4 ) ? ( slice_stream_full ) : ( n403 ) ;
assign n405 =  ( LB2D_shift_x ) >= ( 9'd8 )  ;
assign n406 =  ( LB2D_shift_x ) == ( 9'd0 )  ;
assign n407 =  ( n405 ) | ( n406 )  ;
assign n408 = n127[71:64] ;
assign n409 = LB2D_shift_7[71:64] ;
assign n410 = LB2D_shift_6[71:64] ;
assign n411 = LB2D_shift_5[71:64] ;
assign n412 = LB2D_shift_4[71:64] ;
assign n413 = LB2D_shift_3[71:64] ;
assign n414 = LB2D_shift_2[71:64] ;
assign n415 = LB2D_shift_1[71:64] ;
assign n416 = LB2D_shift_0[71:64] ;
assign n417 =  { ( n415 ) , ( n416 ) }  ;
assign n418 =  { ( n414 ) , ( n417 ) }  ;
assign n419 =  { ( n413 ) , ( n418 ) }  ;
assign n420 =  { ( n412 ) , ( n419 ) }  ;
assign n421 =  { ( n411 ) , ( n420 ) }  ;
assign n422 =  { ( n410 ) , ( n421 ) }  ;
assign n423 =  { ( n409 ) , ( n422 ) }  ;
assign n424 =  { ( n408 ) , ( n423 ) }  ;
assign n425 = n127[63:56] ;
assign n426 = LB2D_shift_7[63:56] ;
assign n427 = LB2D_shift_6[63:56] ;
assign n428 = LB2D_shift_5[63:56] ;
assign n429 = LB2D_shift_4[63:56] ;
assign n430 = LB2D_shift_3[63:56] ;
assign n431 = LB2D_shift_2[63:56] ;
assign n432 = LB2D_shift_1[63:56] ;
assign n433 = LB2D_shift_0[63:56] ;
assign n434 =  { ( n432 ) , ( n433 ) }  ;
assign n435 =  { ( n431 ) , ( n434 ) }  ;
assign n436 =  { ( n430 ) , ( n435 ) }  ;
assign n437 =  { ( n429 ) , ( n436 ) }  ;
assign n438 =  { ( n428 ) , ( n437 ) }  ;
assign n439 =  { ( n427 ) , ( n438 ) }  ;
assign n440 =  { ( n426 ) , ( n439 ) }  ;
assign n441 =  { ( n425 ) , ( n440 ) }  ;
assign n442 = n127[55:48] ;
assign n443 = LB2D_shift_7[55:48] ;
assign n444 = LB2D_shift_6[55:48] ;
assign n445 = LB2D_shift_5[55:48] ;
assign n446 = LB2D_shift_4[55:48] ;
assign n447 = LB2D_shift_3[55:48] ;
assign n448 = LB2D_shift_2[55:48] ;
assign n449 = LB2D_shift_1[55:48] ;
assign n450 = LB2D_shift_0[55:48] ;
assign n451 =  { ( n449 ) , ( n450 ) }  ;
assign n452 =  { ( n448 ) , ( n451 ) }  ;
assign n453 =  { ( n447 ) , ( n452 ) }  ;
assign n454 =  { ( n446 ) , ( n453 ) }  ;
assign n455 =  { ( n445 ) , ( n454 ) }  ;
assign n456 =  { ( n444 ) , ( n455 ) }  ;
assign n457 =  { ( n443 ) , ( n456 ) }  ;
assign n458 =  { ( n442 ) , ( n457 ) }  ;
assign n459 = n127[47:40] ;
assign n460 = LB2D_shift_7[47:40] ;
assign n461 = LB2D_shift_6[47:40] ;
assign n462 = LB2D_shift_5[47:40] ;
assign n463 = LB2D_shift_4[47:40] ;
assign n464 = LB2D_shift_3[47:40] ;
assign n465 = LB2D_shift_2[47:40] ;
assign n466 = LB2D_shift_1[47:40] ;
assign n467 = LB2D_shift_0[47:40] ;
assign n468 =  { ( n466 ) , ( n467 ) }  ;
assign n469 =  { ( n465 ) , ( n468 ) }  ;
assign n470 =  { ( n464 ) , ( n469 ) }  ;
assign n471 =  { ( n463 ) , ( n470 ) }  ;
assign n472 =  { ( n462 ) , ( n471 ) }  ;
assign n473 =  { ( n461 ) , ( n472 ) }  ;
assign n474 =  { ( n460 ) , ( n473 ) }  ;
assign n475 =  { ( n459 ) , ( n474 ) }  ;
assign n476 = n127[39:32] ;
assign n477 = LB2D_shift_7[39:32] ;
assign n478 = LB2D_shift_6[39:32] ;
assign n479 = LB2D_shift_5[39:32] ;
assign n480 = LB2D_shift_4[39:32] ;
assign n481 = LB2D_shift_3[39:32] ;
assign n482 = LB2D_shift_2[39:32] ;
assign n483 = LB2D_shift_1[39:32] ;
assign n484 = LB2D_shift_0[39:32] ;
assign n485 =  { ( n483 ) , ( n484 ) }  ;
assign n486 =  { ( n482 ) , ( n485 ) }  ;
assign n487 =  { ( n481 ) , ( n486 ) }  ;
assign n488 =  { ( n480 ) , ( n487 ) }  ;
assign n489 =  { ( n479 ) , ( n488 ) }  ;
assign n490 =  { ( n478 ) , ( n489 ) }  ;
assign n491 =  { ( n477 ) , ( n490 ) }  ;
assign n492 =  { ( n476 ) , ( n491 ) }  ;
assign n493 = n127[31:24] ;
assign n494 = LB2D_shift_7[31:24] ;
assign n495 = LB2D_shift_6[31:24] ;
assign n496 = LB2D_shift_5[31:24] ;
assign n497 = LB2D_shift_4[31:24] ;
assign n498 = LB2D_shift_3[31:24] ;
assign n499 = LB2D_shift_2[31:24] ;
assign n500 = LB2D_shift_1[31:24] ;
assign n501 = LB2D_shift_0[31:24] ;
assign n502 =  { ( n500 ) , ( n501 ) }  ;
assign n503 =  { ( n499 ) , ( n502 ) }  ;
assign n504 =  { ( n498 ) , ( n503 ) }  ;
assign n505 =  { ( n497 ) , ( n504 ) }  ;
assign n506 =  { ( n496 ) , ( n505 ) }  ;
assign n507 =  { ( n495 ) , ( n506 ) }  ;
assign n508 =  { ( n494 ) , ( n507 ) }  ;
assign n509 =  { ( n493 ) , ( n508 ) }  ;
assign n510 = n127[23:16] ;
assign n511 = LB2D_shift_7[23:16] ;
assign n512 = LB2D_shift_6[23:16] ;
assign n513 = LB2D_shift_5[23:16] ;
assign n514 = LB2D_shift_4[23:16] ;
assign n515 = LB2D_shift_3[23:16] ;
assign n516 = LB2D_shift_2[23:16] ;
assign n517 = LB2D_shift_1[23:16] ;
assign n518 = LB2D_shift_0[23:16] ;
assign n519 =  { ( n517 ) , ( n518 ) }  ;
assign n520 =  { ( n516 ) , ( n519 ) }  ;
assign n521 =  { ( n515 ) , ( n520 ) }  ;
assign n522 =  { ( n514 ) , ( n521 ) }  ;
assign n523 =  { ( n513 ) , ( n522 ) }  ;
assign n524 =  { ( n512 ) , ( n523 ) }  ;
assign n525 =  { ( n511 ) , ( n524 ) }  ;
assign n526 =  { ( n510 ) , ( n525 ) }  ;
assign n527 = n127[15:8] ;
assign n528 = LB2D_shift_7[15:8] ;
assign n529 = LB2D_shift_6[15:8] ;
assign n530 = LB2D_shift_5[15:8] ;
assign n531 = LB2D_shift_4[15:8] ;
assign n532 = LB2D_shift_3[15:8] ;
assign n533 = LB2D_shift_2[15:8] ;
assign n534 = LB2D_shift_1[15:8] ;
assign n535 = LB2D_shift_0[15:8] ;
assign n536 =  { ( n534 ) , ( n535 ) }  ;
assign n537 =  { ( n533 ) , ( n536 ) }  ;
assign n538 =  { ( n532 ) , ( n537 ) }  ;
assign n539 =  { ( n531 ) , ( n538 ) }  ;
assign n540 =  { ( n530 ) , ( n539 ) }  ;
assign n541 =  { ( n529 ) , ( n540 ) }  ;
assign n542 =  { ( n528 ) , ( n541 ) }  ;
assign n543 =  { ( n527 ) , ( n542 ) }  ;
assign n544 = n127[7:0] ;
assign n545 = LB2D_shift_7[7:0] ;
assign n546 = LB2D_shift_6[7:0] ;
assign n547 = LB2D_shift_5[7:0] ;
assign n548 = LB2D_shift_4[7:0] ;
assign n549 = LB2D_shift_3[7:0] ;
assign n550 = LB2D_shift_2[7:0] ;
assign n551 = LB2D_shift_1[7:0] ;
assign n552 = LB2D_shift_0[7:0] ;
assign n553 =  { ( n551 ) , ( n552 ) }  ;
assign n554 =  { ( n550 ) , ( n553 ) }  ;
assign n555 =  { ( n549 ) , ( n554 ) }  ;
assign n556 =  { ( n548 ) , ( n555 ) }  ;
assign n557 =  { ( n547 ) , ( n556 ) }  ;
assign n558 =  { ( n546 ) , ( n557 ) }  ;
assign n559 =  { ( n545 ) , ( n558 ) }  ;
assign n560 =  { ( n544 ) , ( n559 ) }  ;
assign n561 =  { ( n543 ) , ( n560 ) }  ;
assign n562 =  { ( n526 ) , ( n561 ) }  ;
assign n563 =  { ( n509 ) , ( n562 ) }  ;
assign n564 =  { ( n492 ) , ( n563 ) }  ;
assign n565 =  { ( n475 ) , ( n564 ) }  ;
assign n566 =  { ( n458 ) , ( n565 ) }  ;
assign n567 =  { ( n441 ) , ( n566 ) }  ;
assign n568 =  { ( n424 ) , ( n567 ) }  ;
assign n569 =  ( n407 ) ? ( n568 ) : ( stencil_stream_buff_0 ) ;
assign n570 =  ( n34 ) ? ( stencil_stream_buff_0 ) : ( stencil_stream_buff_0 ) ;
assign n571 =  ( n27 ) ? ( stencil_stream_buff_0 ) : ( n570 ) ;
assign n572 =  ( n22 ) ? ( n569 ) : ( n571 ) ;
assign n573 =  ( n13 ) ? ( stencil_stream_buff_0 ) : ( n572 ) ;
assign n574 =  ( n4 ) ? ( stencil_stream_buff_0 ) : ( n573 ) ;
assign n575 =  ( n34 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_1 ) ;
assign n576 =  ( n27 ) ? ( stencil_stream_buff_1 ) : ( n575 ) ;
assign n577 =  ( n22 ) ? ( stencil_stream_buff_0 ) : ( n576 ) ;
assign n578 =  ( n13 ) ? ( stencil_stream_buff_1 ) : ( n577 ) ;
assign n579 =  ( n4 ) ? ( stencil_stream_buff_1 ) : ( n578 ) ;
assign n580 =  ( n154 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n581 = ~ ( n407 ) ;
assign n582 =  ( n581 ) ? ( stencil_stream_empty ) : ( 1'd0 ) ;
assign n583 =  ( n34 ) ? ( stencil_stream_empty ) : ( stencil_stream_empty ) ;
assign n584 =  ( n27 ) ? ( stencil_stream_empty ) : ( n583 ) ;
assign n585 =  ( n22 ) ? ( n582 ) : ( n584 ) ;
assign n586 =  ( n13 ) ? ( n580 ) : ( n585 ) ;
assign n587 =  ( n4 ) ? ( stencil_stream_empty ) : ( n586 ) ;
assign n588 =  ( n9 ) ? ( 1'd0 ) : ( 1'd0 ) ;
assign n589 =  ( stencil_stream_empty ) == ( 1'd1 )  ;
assign n590 =  ( n589 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n591 =  ( n581 ) ? ( stencil_stream_full ) : ( n590 ) ;
assign n592 =  ( n34 ) ? ( stencil_stream_full ) : ( stencil_stream_full ) ;
assign n593 =  ( n27 ) ? ( stencil_stream_full ) : ( n592 ) ;
assign n594 =  ( n22 ) ? ( n591 ) : ( n593 ) ;
assign n595 =  ( n13 ) ? ( n588 ) : ( n594 ) ;
assign n596 =  ( n4 ) ? ( stencil_stream_full ) : ( n595 ) ;
assign n597 = ~ ( n4 ) ;
assign n598 = ~ ( n13 ) ;
assign n599 =  ( n597 ) & ( n598 )  ;
assign n600 = ~ ( n22 ) ;
assign n601 =  ( n599 ) & ( n600 )  ;
assign n602 = ~ ( n27 ) ;
assign n603 =  ( n601 ) & ( n602 )  ;
assign n604 = ~ ( n34 ) ;
assign n605 =  ( n603 ) & ( n604 )  ;
assign n606 =  ( n603 ) & ( n34 )  ;
assign n607 =  ( n601 ) & ( n27 )  ;
assign n608 = ~ ( n298 ) ;
assign n609 =  ( n607 ) & ( n608 )  ;
assign n610 =  ( n607 ) & ( n298 )  ;
assign n611 =  ( n599 ) & ( n22 )  ;
assign n612 =  ( n597 ) & ( n13 )  ;
assign LB2D_proc_0_addr0 = n610 ? (n299) : (0);
assign LB2D_proc_0_data0 = n610 ? (n297) : (LB2D_proc_0[0]);
assign n613 = ~ ( n301 ) ;
assign n614 =  ( n607 ) & ( n613 )  ;
assign n615 =  ( n607 ) & ( n301 )  ;
assign LB2D_proc_1_addr0 = n615 ? (n299) : (0);
assign LB2D_proc_1_data0 = n615 ? (n297) : (LB2D_proc_1[0]);
assign n616 = ~ ( n303 ) ;
assign n617 =  ( n607 ) & ( n616 )  ;
assign n618 =  ( n607 ) & ( n303 )  ;
assign LB2D_proc_2_addr0 = n618 ? (n299) : (0);
assign LB2D_proc_2_data0 = n618 ? (n297) : (LB2D_proc_2[0]);
assign n619 = ~ ( n305 ) ;
assign n620 =  ( n607 ) & ( n619 )  ;
assign n621 =  ( n607 ) & ( n305 )  ;
assign LB2D_proc_3_addr0 = n621 ? (n299) : (0);
assign LB2D_proc_3_data0 = n621 ? (n297) : (LB2D_proc_3[0]);
assign n622 = ~ ( n307 ) ;
assign n623 =  ( n607 ) & ( n622 )  ;
assign n624 =  ( n607 ) & ( n307 )  ;
assign LB2D_proc_4_addr0 = n624 ? (n299) : (0);
assign LB2D_proc_4_data0 = n624 ? (n297) : (LB2D_proc_4[0]);
assign n625 = ~ ( n309 ) ;
assign n626 =  ( n607 ) & ( n625 )  ;
assign n627 =  ( n607 ) & ( n309 )  ;
assign LB2D_proc_5_addr0 = n627 ? (n299) : (0);
assign LB2D_proc_5_data0 = n627 ? (n297) : (LB2D_proc_5[0]);
assign n628 = ~ ( n311 ) ;
assign n629 =  ( n607 ) & ( n628 )  ;
assign n630 =  ( n607 ) & ( n311 )  ;
assign LB2D_proc_6_addr0 = n630 ? (n299) : (0);
assign LB2D_proc_6_data0 = n630 ? (n297) : (LB2D_proc_6[0]);
assign n631 = ~ ( n66 ) ;
assign n632 =  ( n607 ) & ( n631 )  ;
assign n633 =  ( n607 ) & ( n66 )  ;
assign LB2D_proc_7_addr0 = n633 ? (n299) : (0);
assign LB2D_proc_7_data0 = n633 ? (n297) : (LB2D_proc_7[0]);
/*
function [7:0] gb_fun ;
input [647:0] arg0;
    begin
//TODO: Add the specific function HERE.    end
endfunction
*/

always @(posedge clk) begin
   if(rst) begin
       LB1D_buff <= LB1D_buff;
       LB1D_in <= LB1D_in;
       LB1D_it_1 <= LB1D_it_1;
       LB1D_p_cnt <= LB1D_p_cnt;
       LB1D_uIn <= LB1D_uIn;
       LB2D_proc_w <= LB2D_proc_w;
       LB2D_proc_x <= LB2D_proc_x;
       LB2D_proc_y <= LB2D_proc_y;
       LB2D_shift_0 <= LB2D_shift_0;
       LB2D_shift_1 <= LB2D_shift_1;
       LB2D_shift_2 <= LB2D_shift_2;
       LB2D_shift_3 <= LB2D_shift_3;
       LB2D_shift_4 <= LB2D_shift_4;
       LB2D_shift_5 <= LB2D_shift_5;
       LB2D_shift_6 <= LB2D_shift_6;
       LB2D_shift_7 <= LB2D_shift_7;
       LB2D_shift_x <= LB2D_shift_x;
       LB2D_shift_y <= LB2D_shift_y;
       arg_0_TDATA <= arg_0_TDATA;
       arg_0_TVALID <= arg_0_TVALID;
       arg_1_TREADY <= arg_1_TREADY;
       gb_exit_it_1 <= gb_exit_it_1;
       gb_exit_it_2 <= gb_exit_it_2;
       gb_exit_it_3 <= gb_exit_it_3;
       gb_exit_it_4 <= gb_exit_it_4;
       gb_exit_it_5 <= gb_exit_it_5;
       gb_exit_it_6 <= gb_exit_it_6;
       gb_exit_it_7 <= gb_exit_it_7;
       gb_exit_it_8 <= gb_exit_it_8;
       gb_p_cnt <= gb_p_cnt;
       gb_pp_it_1 <= gb_pp_it_1;
       gb_pp_it_2 <= gb_pp_it_2;
       gb_pp_it_3 <= gb_pp_it_3;
       gb_pp_it_4 <= gb_pp_it_4;
       gb_pp_it_5 <= gb_pp_it_5;
       gb_pp_it_6 <= gb_pp_it_6;
       gb_pp_it_7 <= gb_pp_it_7;
       gb_pp_it_8 <= gb_pp_it_8;
       gb_pp_it_9 <= gb_pp_it_9;
       in_stream_buff_0 <= in_stream_buff_0;
       in_stream_buff_1 <= in_stream_buff_1;
       in_stream_empty <= in_stream_empty;
       in_stream_full <= in_stream_full;
       slice_stream_buff_0 <= slice_stream_buff_0;
       slice_stream_buff_1 <= slice_stream_buff_1;
       slice_stream_empty <= slice_stream_empty;
       slice_stream_full <= slice_stream_full;
       stencil_stream_buff_0 <= stencil_stream_buff_0;
       stencil_stream_buff_1 <= stencil_stream_buff_1;
       stencil_stream_empty <= stencil_stream_empty;
       stencil_stream_full <= stencil_stream_full;
   end
   else if(step) begin
       LB1D_buff <= n40;
       LB1D_in <= n46;
       LB1D_it_1 <= n50;
       LB1D_p_cnt <= n58;
       LB1D_uIn <= n64;
       LB2D_proc_w <= n74;
       LB2D_proc_x <= n81;
       LB2D_proc_y <= n90;
       LB2D_shift_0 <= n95;
       LB2D_shift_1 <= n100;
       LB2D_shift_2 <= n105;
       LB2D_shift_3 <= n110;
       LB2D_shift_4 <= n115;
       LB2D_shift_5 <= n120;
       LB2D_shift_6 <= n125;
       LB2D_shift_7 <= n132;
       LB2D_shift_x <= n143;
       LB2D_shift_y <= n153;
       arg_0_TDATA <= n161;
       arg_0_TVALID <= n168;
       arg_1_TREADY <= n177;
       gb_exit_it_1 <= n185;
       gb_exit_it_2 <= n190;
       gb_exit_it_3 <= n195;
       gb_exit_it_4 <= n200;
       gb_exit_it_5 <= n205;
       gb_exit_it_6 <= n210;
       gb_exit_it_7 <= n215;
       gb_exit_it_8 <= n220;
       gb_p_cnt <= n227;
       gb_pp_it_1 <= n232;
       gb_pp_it_2 <= n237;
       gb_pp_it_3 <= n242;
       gb_pp_it_4 <= n247;
       gb_pp_it_5 <= n252;
       gb_pp_it_6 <= n257;
       gb_pp_it_7 <= n262;
       gb_pp_it_8 <= n267;
       gb_pp_it_9 <= n272;
       in_stream_buff_0 <= n277;
       in_stream_buff_1 <= n282;
       in_stream_empty <= n289;
       in_stream_full <= n296;
       slice_stream_buff_0 <= n383;
       slice_stream_buff_1 <= n389;
       slice_stream_empty <= n396;
       slice_stream_full <= n404;
       stencil_stream_buff_0 <= n574;
       stencil_stream_buff_1 <= n579;
       stencil_stream_empty <= n587;
       stencil_stream_full <= n596;
       LB2D_proc_0 [ LB2D_proc_0_addr0 ] <= LB2D_proc_0_data0;
       LB2D_proc_1 [ LB2D_proc_1_addr0 ] <= LB2D_proc_1_data0;
       LB2D_proc_2 [ LB2D_proc_2_addr0 ] <= LB2D_proc_2_data0;
       LB2D_proc_3 [ LB2D_proc_3_addr0 ] <= LB2D_proc_3_data0;
       LB2D_proc_4 [ LB2D_proc_4_addr0 ] <= LB2D_proc_4_data0;
       LB2D_proc_5 [ LB2D_proc_5_addr0 ] <= LB2D_proc_5_data0;
       LB2D_proc_6 [ LB2D_proc_6_addr0 ] <= LB2D_proc_6_data0;
       LB2D_proc_7 [ LB2D_proc_7_addr0 ] <= LB2D_proc_7_data0;
   end
end
endmodule
