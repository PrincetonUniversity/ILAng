module RVCExpander(
  input   clock,
  input   reset,
  input  [31:0] io_in,
  output [31:0] io_out_bits,
  output [4:0] io_out_rd,
  output [4:0] io_out_rs1,
  output [4:0] io_out_rs2,
  output [4:0] io_out_rs3,
  output  io_rvc
);
  wire [1:0] T_12;
  wire  T_14;
  wire [7:0] T_15;
  wire  T_17;
  wire [6:0] T_20;
  wire [3:0] T_21;
  wire [1:0] T_22;
  wire  T_23;
  wire  T_24;
  wire [2:0] T_26;
  wire [5:0] T_27;
  wire [6:0] T_28;
  wire [9:0] T_29;
  wire [2:0] T_33;
  wire [4:0] T_34;
  wire [11:0] T_35;
  wire [14:0] T_36;
  wire [17:0] T_37;
  wire [29:0] T_38;
  wire [4:0] T_46;
  wire [31:0] T_53_bits;
  wire [4:0] T_53_rd;
  wire [4:0] T_53_rs1;
  wire [4:0] T_53_rs2;
  wire [4:0] T_53_rs3;
  wire [1:0] T_59;
  wire [2:0] T_60;
  wire [4:0] T_62;
  wire [7:0] T_63;
  wire [2:0] T_65;
  wire [4:0] T_66;
  wire [11:0] T_72;
  wire [12:0] T_73;
  wire [15:0] T_74;
  wire [27:0] T_75;
  wire [31:0] T_92_bits;
  wire [4:0] T_92_rd;
  wire [4:0] T_92_rs1;
  wire [4:0] T_92_rs2;
  wire [4:0] T_92_rs3;
  wire [3:0] T_103;
  wire [6:0] T_104;
  wire [11:0] T_113;
  wire [11:0] T_114;
  wire [14:0] T_115;
  wire [26:0] T_116;
  wire [31:0] T_133_bits;
  wire [4:0] T_133_rd;
  wire [4:0] T_133_rs1;
  wire [4:0] T_133_rs2;
  wire [4:0] T_133_rs3;
  wire [26:0] T_157;
  wire [31:0] T_174_bits;
  wire [4:0] T_174_rd;
  wire [4:0] T_174_rs1;
  wire [4:0] T_174_rs2;
  wire [4:0] T_174_rs3;
  wire [1:0] T_187;
  wire [4:0] T_202;
  wire [7:0] T_204;
  wire [14:0] T_205;
  wire [6:0] T_206;
  wire [11:0] T_207;
  wire [26:0] T_208;
  wire [31:0] T_225_bits;
  wire [4:0] T_225_rd;
  wire [4:0] T_225_rs1;
  wire [4:0] T_225_rs2;
  wire [4:0] T_225_rs3;
  wire [2:0] T_236;
  wire [4:0] T_249;
  wire [7:0] T_251;
  wire [14:0] T_252;
  wire [7:0] T_253;
  wire [12:0] T_254;
  wire [27:0] T_255;
  wire [31:0] T_272_bits;
  wire [4:0] T_272_rd;
  wire [4:0] T_272_rs1;
  wire [4:0] T_272_rs2;
  wire [4:0] T_272_rs3;
  wire [14:0] T_303;
  wire [26:0] T_306;
  wire [31:0] T_323_bits;
  wire [4:0] T_323_rd;
  wire [4:0] T_323_rs1;
  wire [4:0] T_323_rs2;
  wire [4:0] T_323_rs3;
  wire [14:0] T_354;
  wire [26:0] T_357;
  wire [31:0] T_374_bits;
  wire [4:0] T_374_rd;
  wire [4:0] T_374_rs1;
  wire [4:0] T_374_rs2;
  wire [4:0] T_374_rs3;
  wire  T_380;
  wire [6:0] T_384;
  wire [4:0] T_385;
  wire [11:0] T_386;
  wire [4:0] T_387;
  wire [11:0] T_391;
  wire [16:0] T_392;
  wire [19:0] T_393;
  wire [31:0] T_394;
  wire [31:0] T_407_bits;
  wire [4:0] T_407_rd;
  wire [4:0] T_407_rs1;
  wire [4:0] T_407_rs2;
  wire [4:0] T_407_rs3;
  wire [9:0] T_417;
  wire  T_418;
  wire [1:0] T_419;
  wire  T_421;
  wire  T_422;
  wire  T_423;
  wire [2:0] T_424;
  wire [3:0] T_426;
  wire [1:0] T_427;
  wire [5:0] T_428;
  wire [1:0] T_429;
  wire [10:0] T_430;
  wire [12:0] T_431;
  wire [14:0] T_432;
  wire [20:0] T_433;
  wire  T_434;
  wire [9:0] T_456;
  wire  T_478;
  wire [7:0] T_500;
  wire [12:0] T_503;
  wire [19:0] T_504;
  wire [10:0] T_505;
  wire [11:0] T_506;
  wire [31:0] T_507;
  wire [31:0] T_520_bits;
  wire [4:0] T_520_rd;
  wire [4:0] T_520_rs1;
  wire [4:0] T_520_rs2;
  wire [4:0] T_520_rs3;
  wire [16:0] T_538;
  wire [19:0] T_539;
  wire [31:0] T_540;
  wire [31:0] T_553_bits;
  wire [4:0] T_553_rd;
  wire [4:0] T_553_rs1;
  wire [4:0] T_553_rs2;
  wire [4:0] T_553_rs3;
  wire  T_567;
  wire [6:0] T_570;
  wire [14:0] T_575;
  wire [19:0] T_578;
  wire [31:0] T_579;
  wire [19:0] T_580;
  wire [24:0] T_582;
  wire [31:0] T_583;
  wire [31:0] T_596_bits;
  wire [4:0] T_596_rd;
  wire [4:0] T_596_rs1;
  wire [4:0] T_596_rs2;
  wire [4:0] T_596_rs3;
  wire  T_604;
  wire  T_607;
  wire  T_608;
  wire [6:0] T_620;
  wire [2:0] T_625;
  wire [1:0] T_626;
  wire [1:0] T_631;
  wire [5:0] T_632;
  wire [4:0] T_633;
  wire [5:0] T_634;
  wire [11:0] T_635;
  wire [11:0] T_639;
  wire [16:0] T_640;
  wire [19:0] T_641;
  wire [31:0] T_642;
  wire [31:0] T_655_bits;
  wire [4:0] T_655_rd;
  wire [4:0] T_655_rs1;
  wire [4:0] T_655_rs2;
  wire [4:0] T_655_rs3;
  wire [31:0] T_661_bits;
  wire [4:0] T_661_rd;
  wire [4:0] T_661_rs1;
  wire [4:0] T_661_rs2;
  wire [4:0] T_661_rs3;
  wire [5:0] T_669;
  wire [11:0] T_678;
  wire [10:0] T_679;
  wire [13:0] T_680;
  wire [25:0] T_681;
  wire [30:0] GEN_0;
  wire [30:0] T_698;
  wire [16:0] T_715;
  wire [19:0] T_716;
  wire [31:0] T_717;
  wire [2:0] T_728;
  wire [2:0] T_730;
  wire  T_732;
  wire [2:0] T_734;
  wire  T_736;
  wire  T_740;
  wire [1:0] T_741;
  wire [1:0] T_747;
  wire [2:0] T_756;
  wire [2:0] T_761;
  wire [2:0] T_762;
  wire [2:0] T_763;
  wire  T_766;
  wire [30:0] T_769;
  wire [6:0] T_773;
  wire [11:0] T_783;
  wire [9:0] T_784;
  wire [12:0] T_785;
  wire [24:0] T_786;
  wire [30:0] GEN_1;
  wire [30:0] T_787;
  wire [1:0] T_788;
  wire [1:0] T_790;
  wire  T_792;
  wire  T_796;
  wire [31:0] T_797;
  wire [30:0] T_802;
  wire [31:0] T_803;
  wire [31:0] T_820_bits;
  wire [4:0] T_820_rd;
  wire [4:0] T_820_rs1;
  wire [4:0] T_820_rs2;
  wire [4:0] T_820_rs3;
  wire [12:0] T_916;
  wire [19:0] T_917;
  wire [31:0] T_920;
  wire [31:0] T_935_bits;
  wire [4:0] T_935_rd;
  wire [4:0] T_935_rs1;
  wire [4:0] T_935_rs2;
  wire [4:0] T_935_rs3;
  wire [4:0] T_945;
  wire [3:0] T_951;
  wire [4:0] T_952;
  wire [6:0] T_953;
  wire [7:0] T_954;
  wire [12:0] T_955;
  wire  T_956;
  wire [5:0] T_972;
  wire [3:0] T_993;
  wire  T_1009;
  wire [7:0] T_1011;
  wire [6:0] T_1012;
  wire [14:0] T_1013;
  wire [9:0] T_1014;
  wire [6:0] T_1015;
  wire [16:0] T_1016;
  wire [31:0] T_1017;
  wire [31:0] T_1032_bits;
  wire [4:0] T_1032_rd;
  wire [4:0] T_1032_rs1;
  wire [4:0] T_1032_rs2;
  wire [4:0] T_1032_rs3;
  wire [6:0] T_1109;
  wire [14:0] T_1110;
  wire [31:0] T_1114;
  wire [31:0] T_1127_bits;
  wire [4:0] T_1127_rd;
  wire [4:0] T_1127_rs1;
  wire [4:0] T_1127_rs2;
  wire [4:0] T_1127_rs3;
  wire [10:0] T_1141;
  wire [13:0] T_1142;
  wire [25:0] T_1143;
  wire [31:0] T_1154_bits;
  wire [4:0] T_1154_rd;
  wire [4:0] T_1154_rs1;
  wire [4:0] T_1154_rs2;
  wire [4:0] T_1154_rs3;
  wire [4:0] T_1164;
  wire [3:0] T_1165;
  wire [8:0] T_1166;
  wire [11:0] T_1171;
  wire [13:0] T_1172;
  wire [16:0] T_1173;
  wire [28:0] T_1174;
  wire [31:0] T_1185_bits;
  wire [4:0] T_1185_rd;
  wire [4:0] T_1185_rs1;
  wire [4:0] T_1185_rs2;
  wire [4:0] T_1185_rs3;
  wire [1:0] T_1191;
  wire [2:0] T_1193;
  wire [4:0] T_1195;
  wire [2:0] T_1196;
  wire [7:0] T_1197;
  wire [11:0] T_1202;
  wire [12:0] T_1203;
  wire [15:0] T_1204;
  wire [27:0] T_1205;
  wire [31:0] T_1216_bits;
  wire [4:0] T_1216_rd;
  wire [4:0] T_1216_rs1;
  wire [4:0] T_1216_rs2;
  wire [4:0] T_1216_rs3;
  wire [27:0] T_1236;
  wire [31:0] T_1247_bits;
  wire [4:0] T_1247_rd;
  wire [4:0] T_1247_rs1;
  wire [4:0] T_1247_rs2;
  wire [4:0] T_1247_rs3;
  wire [11:0] T_1258;
  wire [9:0] T_1259;
  wire [12:0] T_1260;
  wire [24:0] T_1261;
  wire [31:0] T_1272_bits;
  wire [4:0] T_1272_rd;
  wire [4:0] T_1272_rs1;
  wire [4:0] T_1272_rs2;
  wire [4:0] T_1272_rs3;
  wire [9:0] T_1284;
  wire [12:0] T_1285;
  wire [24:0] T_1286;
  wire [31:0] T_1297_bits;
  wire [4:0] T_1297_rd;
  wire [4:0] T_1297_rs1;
  wire [4:0] T_1297_rs2;
  wire [4:0] T_1297_rs3;
  wire [24:0] T_1311;
  wire [17:0] T_1312;
  wire [24:0] T_1314;
  wire  T_1317;
  wire [24:0] T_1318;
  wire [31:0] T_1329_bits;
  wire [4:0] T_1329_rd;
  wire [4:0] T_1329_rs1;
  wire [4:0] T_1329_rs2;
  wire [4:0] T_1329_rs3;
  wire  T_1337;
  wire [31:0] T_1338_bits;
  wire [4:0] T_1338_rd;
  wire [4:0] T_1338_rs1;
  wire [4:0] T_1338_rs2;
  wire [4:0] T_1338_rs3;
  wire [24:0] T_1352;
  wire [24:0] T_1355;
  wire [24:0] T_1357;
  wire [24:0] T_1361;
  wire [31:0] T_1372_bits;
  wire [4:0] T_1372_rd;
  wire [4:0] T_1372_rs1;
  wire [4:0] T_1372_rs2;
  wire [4:0] T_1372_rs3;
  wire [31:0] T_1381_bits;
  wire [4:0] T_1381_rd;
  wire [4:0] T_1381_rs1;
  wire [4:0] T_1381_rs2;
  wire [4:0] T_1381_rs3;
  wire [31:0] T_1388_bits;
  wire [4:0] T_1388_rd;
  wire [4:0] T_1388_rs1;
  wire [4:0] T_1388_rs2;
  wire [4:0] T_1388_rs3;
  wire [5:0] T_1397;
  wire [8:0] T_1398;
  wire [3:0] T_1399;
  wire [4:0] T_1408;
  wire [7:0] T_1410;
  wire [14:0] T_1411;
  wire [8:0] T_1412;
  wire [13:0] T_1413;
  wire [28:0] T_1414;
  wire [31:0] T_1425_bits;
  wire [4:0] T_1425_rd;
  wire [4:0] T_1425_rs1;
  wire [4:0] T_1425_rs2;
  wire [4:0] T_1425_rs3;
  wire [1:0] T_1431;
  wire [3:0] T_1432;
  wire [5:0] T_1434;
  wire [7:0] T_1435;
  wire [2:0] T_1436;
  wire [4:0] T_1445;
  wire [7:0] T_1447;
  wire [14:0] T_1448;
  wire [7:0] T_1449;
  wire [12:0] T_1450;
  wire [27:0] T_1451;
  wire [31:0] T_1462_bits;
  wire [4:0] T_1462_rd;
  wire [4:0] T_1462_rs1;
  wire [4:0] T_1462_rs2;
  wire [4:0] T_1462_rs3;
  wire [14:0] T_1485;
  wire [27:0] T_1488;
  wire [31:0] T_1499_bits;
  wire [4:0] T_1499_rd;
  wire [4:0] T_1499_rs1;
  wire [4:0] T_1499_rs2;
  wire [4:0] T_1499_rs3;
  wire [4:0] T_1506;
  wire [4:0] T_1507;
  wire [31:0] T_1515_bits;
  wire [4:0] T_1515_rd;
  wire [4:0] T_1515_rs1;
  wire [4:0] T_1515_rs2;
  wire [4:0] T_1515_rs3;
  wire [31:0] T_1531_bits;
  wire [4:0] T_1531_rd;
  wire [4:0] T_1531_rs1;
  wire [4:0] T_1531_rs2;
  wire [4:0] T_1531_rs3;
  wire [31:0] T_1547_bits;
  wire [4:0] T_1547_rd;
  wire [4:0] T_1547_rs1;
  wire [4:0] T_1547_rs2;
  wire [4:0] T_1547_rs3;
  wire [31:0] T_1563_bits;
  wire [4:0] T_1563_rd;
  wire [4:0] T_1563_rs1;
  wire [4:0] T_1563_rs2;
  wire [4:0] T_1563_rs3;
  wire [31:0] T_1579_bits;
  wire [4:0] T_1579_rd;
  wire [4:0] T_1579_rs1;
  wire [4:0] T_1579_rs2;
  wire [4:0] T_1579_rs3;
  wire [31:0] T_1595_bits;
  wire [4:0] T_1595_rd;
  wire [4:0] T_1595_rs1;
  wire [4:0] T_1595_rs2;
  wire [4:0] T_1595_rs3;
  wire [31:0] T_1611_bits;
  wire [4:0] T_1611_rd;
  wire [4:0] T_1611_rs1;
  wire [4:0] T_1611_rs2;
  wire [4:0] T_1611_rs3;
  wire [31:0] T_1627_bits;
  wire [4:0] T_1627_rd;
  wire [4:0] T_1627_rs1;
  wire [4:0] T_1627_rs2;
  wire [4:0] T_1627_rs3;
  wire [2:0] T_1634;
  wire [4:0] T_1635;
  wire [4:0] T_1637;
  wire  T_1639;
  wire [4:0] T_1641;
  wire  T_1643;
  wire [4:0] T_1645;
  wire  T_1647;
  wire [4:0] T_1649;
  wire  T_1651;
  wire  T_1655;
  wire [31:0] T_1656_bits;
  wire [4:0] T_1656_rd;
  wire [4:0] T_1656_rs1;
  wire [4:0] T_1656_rs2;
  wire [4:0] T_1656_rs3;
  wire [31:0] T_1666_bits;
  wire [4:0] T_1666_rd;
  wire [4:0] T_1666_rs1;
  wire [4:0] T_1666_rs2;
  wire [4:0] T_1666_rs3;
  wire [31:0] T_1672_bits;
  wire [4:0] T_1672_rd;
  wire [4:0] T_1672_rs1;
  wire [4:0] T_1672_rs2;
  wire [4:0] T_1672_rs3;
  wire [31:0] T_1686_bits;
  wire [4:0] T_1686_rd;
  wire [4:0] T_1686_rs1;
  wire [4:0] T_1686_rs2;
  wire [4:0] T_1686_rs3;
  wire [31:0] T_1696_bits;
  wire [4:0] T_1696_rd;
  wire [4:0] T_1696_rs1;
  wire [4:0] T_1696_rs2;
  wire [4:0] T_1696_rs3;
  wire [31:0] T_1702_bits;
  wire [4:0] T_1702_rd;
  wire [4:0] T_1702_rs1;
  wire [4:0] T_1702_rs2;
  wire [4:0] T_1702_rs3;
  wire [31:0] T_1708_bits;
  wire [4:0] T_1708_rd;
  wire [4:0] T_1708_rs1;
  wire [4:0] T_1708_rs2;
  wire [4:0] T_1708_rs3;
  wire [31:0] T_1726_bits;
  wire [4:0] T_1726_rd;
  wire [4:0] T_1726_rs1;
  wire [4:0] T_1726_rs2;
  wire [4:0] T_1726_rs3;
  wire [31:0] T_1736_bits;
  wire [4:0] T_1736_rd;
  wire [4:0] T_1736_rs1;
  wire [4:0] T_1736_rs2;
  wire [4:0] T_1736_rs3;
  wire [31:0] T_1742_bits;
  wire [4:0] T_1742_rd;
  wire [4:0] T_1742_rs1;
  wire [4:0] T_1742_rs2;
  wire [4:0] T_1742_rs3;
  wire [31:0] T_1756_bits;
  wire [4:0] T_1756_rd;
  wire [4:0] T_1756_rs1;
  wire [4:0] T_1756_rs2;
  wire [4:0] T_1756_rs3;
  wire [31:0] T_1766_bits;
  wire [4:0] T_1766_rd;
  wire [4:0] T_1766_rs1;
  wire [4:0] T_1766_rs2;
  wire [4:0] T_1766_rs3;
  wire [31:0] T_1772_bits;
  wire [4:0] T_1772_rd;
  wire [4:0] T_1772_rs1;
  wire [4:0] T_1772_rs2;
  wire [4:0] T_1772_rs3;
  wire [31:0] T_1778_bits;
  wire [4:0] T_1778_rd;
  wire [4:0] T_1778_rs1;
  wire [4:0] T_1778_rs2;
  wire [4:0] T_1778_rs3;
  wire [31:0] T_1784_bits;
  wire [4:0] T_1784_rd;
  wire [4:0] T_1784_rs1;
  wire [4:0] T_1784_rs2;
  wire [4:0] T_1784_rs3;
  wire [31:0] T_1806_bits;
  wire [4:0] T_1806_rd;
  wire [4:0] T_1806_rs1;
  wire [4:0] T_1806_rs2;
  wire [4:0] T_1806_rs3;
  wire [31:0] T_1816_bits;
  wire [4:0] T_1816_rd;
  wire [4:0] T_1816_rs1;
  wire [4:0] T_1816_rs2;
  wire [4:0] T_1816_rs3;
  wire [31:0] T_1822_bits;
  wire [4:0] T_1822_rd;
  wire [4:0] T_1822_rs1;
  wire [4:0] T_1822_rs2;
  wire [4:0] T_1822_rs3;
  wire [31:0] T_1836_bits;
  wire [4:0] T_1836_rd;
  wire [4:0] T_1836_rs1;
  wire [4:0] T_1836_rs2;
  wire [4:0] T_1836_rs3;
  wire [31:0] T_1846_bits;
  wire [4:0] T_1846_rd;
  wire [4:0] T_1846_rs1;
  wire [4:0] T_1846_rs2;
  wire [4:0] T_1846_rs3;
  wire [31:0] T_1852_bits;
  wire [4:0] T_1852_rd;
  wire [4:0] T_1852_rs1;
  wire [4:0] T_1852_rs2;
  wire [4:0] T_1852_rs3;
  wire [31:0] T_1858_bits;
  wire [4:0] T_1858_rd;
  wire [4:0] T_1858_rs1;
  wire [4:0] T_1858_rs2;
  wire [4:0] T_1858_rs3;
  wire [31:0] T_1876_bits;
  wire [4:0] T_1876_rd;
  wire [4:0] T_1876_rs1;
  wire [4:0] T_1876_rs2;
  wire [4:0] T_1876_rs3;
  wire [31:0] T_1886_bits;
  wire [4:0] T_1886_rd;
  wire [4:0] T_1886_rs1;
  wire [4:0] T_1886_rs2;
  wire [4:0] T_1886_rs3;
  wire [31:0] T_1892_bits;
  wire [4:0] T_1892_rd;
  wire [4:0] T_1892_rs1;
  wire [4:0] T_1892_rs2;
  wire [4:0] T_1892_rs3;
  wire [31:0] T_1906_bits;
  wire [4:0] T_1906_rd;
  wire [4:0] T_1906_rs1;
  wire [4:0] T_1906_rs2;
  wire [4:0] T_1906_rs3;
  wire [31:0] T_1916_bits;
  wire [4:0] T_1916_rd;
  wire [4:0] T_1916_rs1;
  wire [4:0] T_1916_rs2;
  wire [4:0] T_1916_rs3;
  wire [31:0] T_1922_bits;
  wire [4:0] T_1922_rd;
  wire [4:0] T_1922_rs1;
  wire [4:0] T_1922_rs2;
  wire [4:0] T_1922_rs3;
  wire [31:0] T_1928_bits;
  wire [4:0] T_1928_rd;
  wire [4:0] T_1928_rs1;
  wire [4:0] T_1928_rs2;
  wire [4:0] T_1928_rs3;
  wire [31:0] T_1934_bits;
  wire [4:0] T_1934_rd;
  wire [4:0] T_1934_rs1;
  wire [4:0] T_1934_rs2;
  wire [4:0] T_1934_rs3;
  wire [31:0] T_1940_bits;
  wire [4:0] T_1940_rd;
  wire [4:0] T_1940_rs1;
  wire [4:0] T_1940_rs2;
  wire [4:0] T_1940_rs3;
  assign io_out_bits = T_1940_bits;
  assign io_out_rd = T_1940_rd;
  assign io_out_rs1 = T_1940_rs1;
  assign io_out_rs2 = T_1940_rs2;
  assign io_out_rs3 = T_1940_rs3;
  assign io_rvc = T_14;
  assign T_12 = io_in[1:0];
  assign T_14 = T_12 != 2'h3;
  assign T_15 = io_in[12:5];
  assign T_17 = T_15 != 8'h0;
  assign T_20 = T_17 ? 7'h13 : 7'h1f;
  assign T_21 = io_in[10:7];
  assign T_22 = io_in[12:11];
  assign T_23 = io_in[5];
  assign T_24 = io_in[6];
  assign T_26 = {T_24,2'h0};
  assign T_27 = {T_21,T_22};
  assign T_28 = {T_27,T_23};
  assign T_29 = {T_28,T_26};
  assign T_33 = io_in[4:2];
  assign T_34 = {2'h1,T_33};
  assign T_35 = {T_34,T_20};
  assign T_36 = {T_29,5'h2};
  assign T_37 = {T_36,3'h0};
  assign T_38 = {T_37,T_35};
  assign T_46 = io_in[31:27];
  assign T_53_bits = {{2'd0}, T_38};
  assign T_53_rd = T_34;
  assign T_53_rs1 = 5'h2;
  assign T_53_rs2 = T_34;
  assign T_53_rs3 = T_46;
  assign T_59 = io_in[6:5];
  assign T_60 = io_in[12:10];
  assign T_62 = {T_59,T_60};
  assign T_63 = {T_62,3'h0};
  assign T_65 = io_in[9:7];
  assign T_66 = {2'h1,T_65};
  assign T_72 = {T_34,7'h7};
  assign T_73 = {T_63,T_66};
  assign T_74 = {T_73,3'h3};
  assign T_75 = {T_74,T_72};
  assign T_92_bits = {{4'd0}, T_75};
  assign T_92_rd = T_34;
  assign T_92_rs1 = T_66;
  assign T_92_rs2 = T_34;
  assign T_92_rs3 = T_46;
  assign T_103 = {T_23,T_60};
  assign T_104 = {T_103,T_26};
  assign T_113 = {T_34,7'h3};
  assign T_114 = {T_104,T_66};
  assign T_115 = {T_114,3'h2};
  assign T_116 = {T_115,T_113};
  assign T_133_bits = {{5'd0}, T_116};
  assign T_133_rd = T_34;
  assign T_133_rs1 = T_66;
  assign T_133_rs2 = T_34;
  assign T_133_rs3 = T_46;
  assign T_157 = {T_115,T_72};
  assign T_174_bits = {{5'd0}, T_157};
  assign T_174_rd = T_34;
  assign T_174_rs1 = T_66;
  assign T_174_rs2 = T_34;
  assign T_174_rs3 = T_46;
  assign T_187 = T_104[6:5];
  assign T_202 = T_104[4:0];
  assign T_204 = {3'h2,T_202};
  assign T_205 = {T_204,7'h2f};
  assign T_206 = {T_187,T_34};
  assign T_207 = {T_206,T_66};
  assign T_208 = {T_207,T_205};
  assign T_225_bits = {{5'd0}, T_208};
  assign T_225_rd = T_34;
  assign T_225_rs1 = T_66;
  assign T_225_rs2 = T_34;
  assign T_225_rs3 = T_46;
  assign T_236 = T_63[7:5];
  assign T_249 = T_63[4:0];
  assign T_251 = {3'h3,T_249};
  assign T_252 = {T_251,7'h27};
  assign T_253 = {T_236,T_34};
  assign T_254 = {T_253,T_66};
  assign T_255 = {T_254,T_252};
  assign T_272_bits = {{4'd0}, T_255};
  assign T_272_rd = T_34;
  assign T_272_rs1 = T_66;
  assign T_272_rs2 = T_34;
  assign T_272_rs3 = T_46;
  assign T_303 = {T_204,7'h23};
  assign T_306 = {T_207,T_303};
  assign T_323_bits = {{5'd0}, T_306};
  assign T_323_rd = T_34;
  assign T_323_rs1 = T_66;
  assign T_323_rs2 = T_34;
  assign T_323_rs3 = T_46;
  assign T_354 = {T_204,7'h27};
  assign T_357 = {T_207,T_354};
  assign T_374_bits = {{5'd0}, T_357};
  assign T_374_rd = T_34;
  assign T_374_rs1 = T_66;
  assign T_374_rs2 = T_34;
  assign T_374_rs3 = T_46;
  assign T_380 = io_in[12];
  assign T_384 = T_380 ? 7'h7f : 7'h0;
  assign T_385 = io_in[6:2];
  assign T_386 = {T_384,T_385};
  assign T_387 = io_in[11:7];
  assign T_391 = {T_387,7'h13};
  assign T_392 = {T_386,T_387};
  assign T_393 = {T_392,3'h0};
  assign T_394 = {T_393,T_391};
  assign T_407_bits = T_394;
  assign T_407_rd = T_387;
  assign T_407_rs1 = T_387;
  assign T_407_rs2 = T_34;
  assign T_407_rs3 = T_46;
  assign T_417 = T_380 ? 10'h3ff : 10'h0;
  assign T_418 = io_in[8];
  assign T_419 = io_in[10:9];
  assign T_421 = io_in[7];
  assign T_422 = io_in[2];
  assign T_423 = io_in[11];
  assign T_424 = io_in[5:3];
  assign T_426 = {T_424,1'h0};
  assign T_427 = {T_422,T_423};
  assign T_428 = {T_427,T_426};
  assign T_429 = {T_24,T_421};
  assign T_430 = {T_417,T_418};
  assign T_431 = {T_430,T_419};
  assign T_432 = {T_431,T_429};
  assign T_433 = {T_432,T_428};
  assign T_434 = T_433[20];
  assign T_456 = T_433[10:1];
  assign T_478 = T_433[11];
  assign T_500 = T_433[19:12];
  assign T_503 = {T_500,5'h1};
  assign T_504 = {T_503,7'h6f};
  assign T_505 = {T_434,T_456};
  assign T_506 = {T_505,T_478};
  assign T_507 = {T_506,T_504};
  assign T_520_bits = T_507;
  assign T_520_rd = 5'h1;
  assign T_520_rs1 = T_387;
  assign T_520_rs2 = T_34;
  assign T_520_rs3 = T_46;
  assign T_538 = {T_386,5'h0};
  assign T_539 = {T_538,3'h0};
  assign T_540 = {T_539,T_391};
  assign T_553_bits = T_540;
  assign T_553_rd = T_387;
  assign T_553_rs1 = 5'h0;
  assign T_553_rs2 = T_34;
  assign T_553_rs3 = T_46;
  assign T_567 = T_386 != 12'h0;
  assign T_570 = T_567 ? 7'h37 : 7'h3f;
  assign T_575 = T_380 ? 15'h7fff : 15'h0;
  assign T_578 = {T_575,T_385};
  assign T_579 = {T_578,12'h0};
  assign T_580 = T_579[31:12];
  assign T_582 = {T_580,T_387};
  assign T_583 = {T_582,T_570};
  assign T_596_bits = T_583;
  assign T_596_rd = T_387;
  assign T_596_rs1 = T_387;
  assign T_596_rs2 = T_34;
  assign T_596_rs3 = T_46;
  assign T_604 = T_387 == 5'h0;
  assign T_607 = T_387 == 5'h2;
  assign T_608 = T_604 | T_607;
  assign T_620 = T_567 ? 7'h13 : 7'h1f;
  assign T_625 = T_380 ? 3'h7 : 3'h0;
  assign T_626 = io_in[4:3];
  assign T_631 = {T_422,T_24};
  assign T_632 = {T_631,4'h0};
  assign T_633 = {T_625,T_626};
  assign T_634 = {T_633,T_23};
  assign T_635 = {T_634,T_632};
  assign T_639 = {T_387,T_620};
  assign T_640 = {T_635,T_387};
  assign T_641 = {T_640,3'h0};
  assign T_642 = {T_641,T_639};
  assign T_655_bits = T_642;
  assign T_655_rd = T_387;
  assign T_655_rs1 = T_387;
  assign T_655_rs2 = T_34;
  assign T_655_rs3 = T_46;
  assign T_661_bits = T_608 ? T_655_bits : T_596_bits;
  assign T_661_rd = T_608 ? T_655_rd : T_596_rd;
  assign T_661_rs1 = T_608 ? T_655_rs1 : T_596_rs1;
  assign T_661_rs2 = T_608 ? T_655_rs2 : T_596_rs2;
  assign T_661_rs3 = T_608 ? T_655_rs3 : T_596_rs3;
  assign T_669 = {T_380,T_385};
  assign T_678 = {T_66,7'h13};
  assign T_679 = {T_669,T_66};
  assign T_680 = {T_679,3'h5};
  assign T_681 = {T_680,T_678};
  assign GEN_0 = {{5'd0}, T_681};
  assign T_698 = GEN_0 | 31'h40000000;
  assign T_715 = {T_386,T_66};
  assign T_716 = {T_715,3'h7};
  assign T_717 = {T_716,T_678};
  assign T_728 = {T_380,T_59};
  assign T_730 = T_728 & 3'h3;
  assign T_732 = T_728 >= 3'h4;
  assign T_734 = T_730 & 3'h1;
  assign T_736 = T_730 >= 3'h2;
  assign T_740 = T_734 >= 3'h1;
  assign T_741 = T_740 ? 2'h3 : 2'h2;
  assign T_747 = T_736 ? T_741 : 2'h0;
  assign T_756 = T_740 ? 3'h7 : 3'h6;
  assign T_761 = T_740 ? 3'h4 : 3'h0;
  assign T_762 = T_736 ? T_756 : T_761;
  assign T_763 = T_732 ? {{1'd0}, T_747} : T_762;
  assign T_766 = T_59 == 2'h0;
  assign T_769 = T_766 ? 31'h40000000 : 31'h0;
  assign T_773 = T_380 ? 7'h3b : 7'h33;
  assign T_783 = {T_66,T_773};
  assign T_784 = {T_34,T_66};
  assign T_785 = {T_784,T_763};
  assign T_786 = {T_785,T_783};
  assign GEN_1 = {{6'd0}, T_786};
  assign T_787 = GEN_1 | T_769;
  assign T_788 = io_in[11:10];
  assign T_790 = T_788 & 2'h1;
  assign T_792 = T_788 >= 2'h2;
  assign T_796 = T_790 >= 2'h1;
  assign T_797 = T_796 ? {{1'd0}, T_787} : T_717;
  assign T_802 = T_796 ? T_698 : {{5'd0}, T_681};
  assign T_803 = T_792 ? T_797 : {{1'd0}, T_802};
  assign T_820_bits = T_803;
  assign T_820_rd = T_66;
  assign T_820_rs1 = T_66;
  assign T_820_rs2 = T_34;
  assign T_820_rs3 = T_46;
  assign T_916 = {T_500,5'h0};
  assign T_917 = {T_916,7'h6f};
  assign T_920 = {T_506,T_917};
  assign T_935_bits = T_920;
  assign T_935_rd = 5'h0;
  assign T_935_rs1 = T_66;
  assign T_935_rs2 = T_34;
  assign T_935_rs3 = T_46;
  assign T_945 = T_380 ? 5'h1f : 5'h0;
  assign T_951 = {T_788,T_626};
  assign T_952 = {T_951,1'h0};
  assign T_953 = {T_945,T_59};
  assign T_954 = {T_953,T_422};
  assign T_955 = {T_954,T_952};
  assign T_956 = T_955[12];
  assign T_972 = T_955[10:5];
  assign T_993 = T_955[4:1];
  assign T_1009 = T_955[11];
  assign T_1011 = {T_1009,7'h63};
  assign T_1012 = {3'h0,T_993};
  assign T_1013 = {T_1012,T_1011};
  assign T_1014 = {5'h0,T_66};
  assign T_1015 = {T_956,T_972};
  assign T_1016 = {T_1015,T_1014};
  assign T_1017 = {T_1016,T_1013};
  assign T_1032_bits = T_1017;
  assign T_1032_rd = T_66;
  assign T_1032_rs1 = T_66;
  assign T_1032_rs2 = 5'h0;
  assign T_1032_rs3 = T_46;
  assign T_1109 = {3'h1,T_993};
  assign T_1110 = {T_1109,T_1011};
  assign T_1114 = {T_1016,T_1110};
  assign T_1127_bits = T_1114;
  assign T_1127_rd = 5'h0;
  assign T_1127_rs1 = T_66;
  assign T_1127_rs2 = 5'h0;
  assign T_1127_rs3 = T_46;
  assign T_1141 = {T_669,T_387};
  assign T_1142 = {T_1141,3'h1};
  assign T_1143 = {T_1142,T_391};
  assign T_1154_bits = {{6'd0}, T_1143};
  assign T_1154_rd = T_387;
  assign T_1154_rs1 = T_387;
  assign T_1154_rs2 = T_385;
  assign T_1154_rs3 = T_46;
  assign T_1164 = {T_59,3'h0};
  assign T_1165 = {T_33,T_380};
  assign T_1166 = {T_1165,T_1164};
  assign T_1171 = {T_387,7'h7};
  assign T_1172 = {T_1166,5'h2};
  assign T_1173 = {T_1172,3'h3};
  assign T_1174 = {T_1173,T_1171};
  assign T_1185_bits = {{3'd0}, T_1174};
  assign T_1185_rd = T_387;
  assign T_1185_rs1 = 5'h2;
  assign T_1185_rs2 = T_385;
  assign T_1185_rs3 = T_46;
  assign T_1191 = io_in[3:2];
  assign T_1193 = io_in[6:4];
  assign T_1195 = {T_1193,2'h0};
  assign T_1196 = {T_1191,T_380};
  assign T_1197 = {T_1196,T_1195};
  assign T_1202 = {T_387,7'h3};
  assign T_1203 = {T_1197,5'h2};
  assign T_1204 = {T_1203,3'h2};
  assign T_1205 = {T_1204,T_1202};
  assign T_1216_bits = {{4'd0}, T_1205};
  assign T_1216_rd = T_387;
  assign T_1216_rs1 = 5'h2;
  assign T_1216_rs2 = T_385;
  assign T_1216_rs3 = T_46;
  assign T_1236 = {T_1204,T_1171};
  assign T_1247_bits = {{4'd0}, T_1236};
  assign T_1247_rd = T_387;
  assign T_1247_rs1 = 5'h2;
  assign T_1247_rs2 = T_385;
  assign T_1247_rs3 = T_46;
  assign T_1258 = {T_387,7'h33};
  assign T_1259 = {T_385,5'h0};
  assign T_1260 = {T_1259,3'h0};
  assign T_1261 = {T_1260,T_1258};
  assign T_1272_bits = {{7'd0}, T_1261};
  assign T_1272_rd = T_387;
  assign T_1272_rs1 = 5'h0;
  assign T_1272_rs2 = T_385;
  assign T_1272_rs3 = T_46;
  assign T_1284 = {T_385,T_387};
  assign T_1285 = {T_1284,3'h0};
  assign T_1286 = {T_1285,T_1258};
  assign T_1297_bits = {{7'd0}, T_1286};
  assign T_1297_rd = T_387;
  assign T_1297_rs1 = T_387;
  assign T_1297_rs2 = T_385;
  assign T_1297_rs3 = T_46;
  assign T_1311 = {T_1285,12'h67};
  assign T_1312 = T_1311[24:7];
  assign T_1314 = {T_1312,7'h1f};
  assign T_1317 = T_387 != 5'h0;
  assign T_1318 = T_1317 ? T_1311 : T_1314;
  assign T_1329_bits = {{7'd0}, T_1318};
  assign T_1329_rd = 5'h0;
  assign T_1329_rs1 = T_387;
  assign T_1329_rs2 = T_385;
  assign T_1329_rs3 = T_46;
  assign T_1337 = T_385 != 5'h0;
  assign T_1338_bits = T_1337 ? T_1272_bits : T_1329_bits;
  assign T_1338_rd = T_1337 ? T_1272_rd : T_1329_rd;
  assign T_1338_rs1 = T_1337 ? T_1272_rs1 : T_1329_rs1;
  assign T_1338_rs2 = T_1337 ? T_1272_rs2 : T_1329_rs2;
  assign T_1338_rs3 = T_1337 ? T_1272_rs3 : T_1329_rs3;
  assign T_1352 = {T_1285,12'he7};
  assign T_1355 = {T_1312,7'h73};
  assign T_1357 = T_1355 | 25'h100000;
  assign T_1361 = T_1317 ? T_1352 : T_1357;
  assign T_1372_bits = {{7'd0}, T_1361};
  assign T_1372_rd = 5'h1;
  assign T_1372_rs1 = T_387;
  assign T_1372_rs2 = T_385;
  assign T_1372_rs3 = T_46;
  assign T_1381_bits = T_1337 ? T_1297_bits : T_1372_bits;
  assign T_1381_rd = T_1337 ? T_1297_rd : T_1372_rd;
  assign T_1381_rs1 = T_1337 ? T_1297_rs1 : T_1372_rs1;
  assign T_1381_rs2 = T_1337 ? T_1297_rs2 : T_1372_rs2;
  assign T_1381_rs3 = T_1337 ? T_1297_rs3 : T_1372_rs3;
  assign T_1388_bits = T_380 ? T_1381_bits : T_1338_bits;
  assign T_1388_rd = T_380 ? T_1381_rd : T_1338_rd;
  assign T_1388_rs1 = T_380 ? T_1381_rs1 : T_1338_rs1;
  assign T_1388_rs2 = T_380 ? T_1381_rs2 : T_1338_rs2;
  assign T_1388_rs3 = T_380 ? T_1381_rs3 : T_1338_rs3;
  assign T_1397 = {T_65,T_60};
  assign T_1398 = {T_1397,3'h0};
  assign T_1399 = T_1398[8:5];
  assign T_1408 = T_1398[4:0];
  assign T_1410 = {3'h3,T_1408};
  assign T_1411 = {T_1410,7'h27};
  assign T_1412 = {T_1399,T_385};
  assign T_1413 = {T_1412,5'h2};
  assign T_1414 = {T_1413,T_1411};
  assign T_1425_bits = {{3'd0}, T_1414};
  assign T_1425_rd = T_387;
  assign T_1425_rs1 = 5'h2;
  assign T_1425_rs2 = T_385;
  assign T_1425_rs3 = T_46;
  assign T_1431 = io_in[8:7];
  assign T_1432 = io_in[12:9];
  assign T_1434 = {T_1431,T_1432};
  assign T_1435 = {T_1434,2'h0};
  assign T_1436 = T_1435[7:5];
  assign T_1445 = T_1435[4:0];
  assign T_1447 = {3'h2,T_1445};
  assign T_1448 = {T_1447,7'h23};
  assign T_1449 = {T_1436,T_385};
  assign T_1450 = {T_1449,5'h2};
  assign T_1451 = {T_1450,T_1448};
  assign T_1462_bits = {{4'd0}, T_1451};
  assign T_1462_rd = T_387;
  assign T_1462_rs1 = 5'h2;
  assign T_1462_rs2 = T_385;
  assign T_1462_rs3 = T_46;
  assign T_1485 = {T_1447,7'h27};
  assign T_1488 = {T_1450,T_1485};
  assign T_1499_bits = {{4'd0}, T_1488};
  assign T_1499_rd = T_387;
  assign T_1499_rs1 = 5'h2;
  assign T_1499_rs2 = T_385;
  assign T_1499_rs3 = T_46;
  assign T_1506 = io_in[19:15];
  assign T_1507 = io_in[24:20];
  assign T_1515_bits = io_in;
  assign T_1515_rd = T_387;
  assign T_1515_rs1 = T_1506;
  assign T_1515_rs2 = T_1507;
  assign T_1515_rs3 = T_46;
  assign T_1531_bits = io_in;
  assign T_1531_rd = T_387;
  assign T_1531_rs1 = T_1506;
  assign T_1531_rs2 = T_1507;
  assign T_1531_rs3 = T_46;
  assign T_1547_bits = io_in;
  assign T_1547_rd = T_387;
  assign T_1547_rs1 = T_1506;
  assign T_1547_rs2 = T_1507;
  assign T_1547_rs3 = T_46;
  assign T_1563_bits = io_in;
  assign T_1563_rd = T_387;
  assign T_1563_rs1 = T_1506;
  assign T_1563_rs2 = T_1507;
  assign T_1563_rs3 = T_46;
  assign T_1579_bits = io_in;
  assign T_1579_rd = T_387;
  assign T_1579_rs1 = T_1506;
  assign T_1579_rs2 = T_1507;
  assign T_1579_rs3 = T_46;
  assign T_1595_bits = io_in;
  assign T_1595_rd = T_387;
  assign T_1595_rs1 = T_1506;
  assign T_1595_rs2 = T_1507;
  assign T_1595_rs3 = T_46;
  assign T_1611_bits = io_in;
  assign T_1611_rd = T_387;
  assign T_1611_rs1 = T_1506;
  assign T_1611_rs2 = T_1507;
  assign T_1611_rs3 = T_46;
  assign T_1627_bits = io_in;
  assign T_1627_rd = T_387;
  assign T_1627_rs1 = T_1506;
  assign T_1627_rs2 = T_1507;
  assign T_1627_rs3 = T_46;
  assign T_1634 = io_in[15:13];
  assign T_1635 = {T_12,T_1634};
  assign T_1637 = T_1635 & 5'hf;
  assign T_1639 = T_1635 >= 5'h10;
  assign T_1641 = T_1637 & 5'h7;
  assign T_1643 = T_1637 >= 5'h8;
  assign T_1645 = T_1641 & 5'h3;
  assign T_1647 = T_1641 >= 5'h4;
  assign T_1649 = T_1645 & 5'h1;
  assign T_1651 = T_1645 >= 5'h2;
  assign T_1655 = T_1649 >= 5'h1;
  assign T_1656_bits = T_1655 ? T_1627_bits : T_1611_bits;
  assign T_1656_rd = T_1655 ? T_1627_rd : T_1611_rd;
  assign T_1656_rs1 = T_1655 ? T_1627_rs1 : T_1611_rs1;
  assign T_1656_rs2 = T_1655 ? T_1627_rs2 : T_1611_rs2;
  assign T_1656_rs3 = T_1655 ? T_1627_rs3 : T_1611_rs3;
  assign T_1666_bits = T_1655 ? T_1595_bits : T_1579_bits;
  assign T_1666_rd = T_1655 ? T_1595_rd : T_1579_rd;
  assign T_1666_rs1 = T_1655 ? T_1595_rs1 : T_1579_rs1;
  assign T_1666_rs2 = T_1655 ? T_1595_rs2 : T_1579_rs2;
  assign T_1666_rs3 = T_1655 ? T_1595_rs3 : T_1579_rs3;
  assign T_1672_bits = T_1651 ? T_1656_bits : T_1666_bits;
  assign T_1672_rd = T_1651 ? T_1656_rd : T_1666_rd;
  assign T_1672_rs1 = T_1651 ? T_1656_rs1 : T_1666_rs1;
  assign T_1672_rs2 = T_1651 ? T_1656_rs2 : T_1666_rs2;
  assign T_1672_rs3 = T_1651 ? T_1656_rs3 : T_1666_rs3;
  assign T_1686_bits = T_1655 ? T_1563_bits : T_1547_bits;
  assign T_1686_rd = T_1655 ? T_1563_rd : T_1547_rd;
  assign T_1686_rs1 = T_1655 ? T_1563_rs1 : T_1547_rs1;
  assign T_1686_rs2 = T_1655 ? T_1563_rs2 : T_1547_rs2;
  assign T_1686_rs3 = T_1655 ? T_1563_rs3 : T_1547_rs3;
  assign T_1696_bits = T_1655 ? T_1531_bits : T_1515_bits;
  assign T_1696_rd = T_1655 ? T_1531_rd : T_1515_rd;
  assign T_1696_rs1 = T_1655 ? T_1531_rs1 : T_1515_rs1;
  assign T_1696_rs2 = T_1655 ? T_1531_rs2 : T_1515_rs2;
  assign T_1696_rs3 = T_1655 ? T_1531_rs3 : T_1515_rs3;
  assign T_1702_bits = T_1651 ? T_1686_bits : T_1696_bits;
  assign T_1702_rd = T_1651 ? T_1686_rd : T_1696_rd;
  assign T_1702_rs1 = T_1651 ? T_1686_rs1 : T_1696_rs1;
  assign T_1702_rs2 = T_1651 ? T_1686_rs2 : T_1696_rs2;
  assign T_1702_rs3 = T_1651 ? T_1686_rs3 : T_1696_rs3;
  assign T_1708_bits = T_1647 ? T_1672_bits : T_1702_bits;
  assign T_1708_rd = T_1647 ? T_1672_rd : T_1702_rd;
  assign T_1708_rs1 = T_1647 ? T_1672_rs1 : T_1702_rs1;
  assign T_1708_rs2 = T_1647 ? T_1672_rs2 : T_1702_rs2;
  assign T_1708_rs3 = T_1647 ? T_1672_rs3 : T_1702_rs3;
  assign T_1726_bits = T_1655 ? T_1499_bits : T_1462_bits;
  assign T_1726_rd = T_1655 ? T_1499_rd : T_1462_rd;
  assign T_1726_rs1 = T_1655 ? T_1499_rs1 : T_1462_rs1;
  assign T_1726_rs2 = T_1655 ? T_1499_rs2 : T_1462_rs2;
  assign T_1726_rs3 = T_1655 ? T_1499_rs3 : T_1462_rs3;
  assign T_1736_bits = T_1655 ? T_1425_bits : T_1388_bits;
  assign T_1736_rd = T_1655 ? T_1425_rd : T_1388_rd;
  assign T_1736_rs1 = T_1655 ? T_1425_rs1 : T_1388_rs1;
  assign T_1736_rs2 = T_1655 ? T_1425_rs2 : T_1388_rs2;
  assign T_1736_rs3 = T_1655 ? T_1425_rs3 : T_1388_rs3;
  assign T_1742_bits = T_1651 ? T_1726_bits : T_1736_bits;
  assign T_1742_rd = T_1651 ? T_1726_rd : T_1736_rd;
  assign T_1742_rs1 = T_1651 ? T_1726_rs1 : T_1736_rs1;
  assign T_1742_rs2 = T_1651 ? T_1726_rs2 : T_1736_rs2;
  assign T_1742_rs3 = T_1651 ? T_1726_rs3 : T_1736_rs3;
  assign T_1756_bits = T_1655 ? T_1247_bits : T_1216_bits;
  assign T_1756_rd = T_1655 ? T_1247_rd : T_1216_rd;
  assign T_1756_rs1 = T_1655 ? T_1247_rs1 : T_1216_rs1;
  assign T_1756_rs2 = T_1655 ? T_1247_rs2 : T_1216_rs2;
  assign T_1756_rs3 = T_1655 ? T_1247_rs3 : T_1216_rs3;
  assign T_1766_bits = T_1655 ? T_1185_bits : T_1154_bits;
  assign T_1766_rd = T_1655 ? T_1185_rd : T_1154_rd;
  assign T_1766_rs1 = T_1655 ? T_1185_rs1 : T_1154_rs1;
  assign T_1766_rs2 = T_1655 ? T_1185_rs2 : T_1154_rs2;
  assign T_1766_rs3 = T_1655 ? T_1185_rs3 : T_1154_rs3;
  assign T_1772_bits = T_1651 ? T_1756_bits : T_1766_bits;
  assign T_1772_rd = T_1651 ? T_1756_rd : T_1766_rd;
  assign T_1772_rs1 = T_1651 ? T_1756_rs1 : T_1766_rs1;
  assign T_1772_rs2 = T_1651 ? T_1756_rs2 : T_1766_rs2;
  assign T_1772_rs3 = T_1651 ? T_1756_rs3 : T_1766_rs3;
  assign T_1778_bits = T_1647 ? T_1742_bits : T_1772_bits;
  assign T_1778_rd = T_1647 ? T_1742_rd : T_1772_rd;
  assign T_1778_rs1 = T_1647 ? T_1742_rs1 : T_1772_rs1;
  assign T_1778_rs2 = T_1647 ? T_1742_rs2 : T_1772_rs2;
  assign T_1778_rs3 = T_1647 ? T_1742_rs3 : T_1772_rs3;
  assign T_1784_bits = T_1643 ? T_1708_bits : T_1778_bits;
  assign T_1784_rd = T_1643 ? T_1708_rd : T_1778_rd;
  assign T_1784_rs1 = T_1643 ? T_1708_rs1 : T_1778_rs1;
  assign T_1784_rs2 = T_1643 ? T_1708_rs2 : T_1778_rs2;
  assign T_1784_rs3 = T_1643 ? T_1708_rs3 : T_1778_rs3;
  assign T_1806_bits = T_1655 ? T_1127_bits : T_1032_bits;
  assign T_1806_rd = T_1655 ? T_1127_rd : T_1032_rd;
  assign T_1806_rs1 = T_1655 ? T_1127_rs1 : T_1032_rs1;
  assign T_1806_rs2 = T_1655 ? T_1127_rs2 : T_1032_rs2;
  assign T_1806_rs3 = T_1655 ? T_1127_rs3 : T_1032_rs3;
  assign T_1816_bits = T_1655 ? T_935_bits : T_820_bits;
  assign T_1816_rd = T_1655 ? T_935_rd : T_820_rd;
  assign T_1816_rs1 = T_1655 ? T_935_rs1 : T_820_rs1;
  assign T_1816_rs2 = T_1655 ? T_935_rs2 : T_820_rs2;
  assign T_1816_rs3 = T_1655 ? T_935_rs3 : T_820_rs3;
  assign T_1822_bits = T_1651 ? T_1806_bits : T_1816_bits;
  assign T_1822_rd = T_1651 ? T_1806_rd : T_1816_rd;
  assign T_1822_rs1 = T_1651 ? T_1806_rs1 : T_1816_rs1;
  assign T_1822_rs2 = T_1651 ? T_1806_rs2 : T_1816_rs2;
  assign T_1822_rs3 = T_1651 ? T_1806_rs3 : T_1816_rs3;
  assign T_1836_bits = T_1655 ? T_661_bits : T_553_bits;
  assign T_1836_rd = T_1655 ? T_661_rd : T_553_rd;
  assign T_1836_rs1 = T_1655 ? T_661_rs1 : T_553_rs1;
  assign T_1836_rs2 = T_1655 ? T_661_rs2 : T_553_rs2;
  assign T_1836_rs3 = T_1655 ? T_661_rs3 : T_553_rs3;
  assign T_1846_bits = T_1655 ? T_520_bits : T_407_bits;
  assign T_1846_rd = T_1655 ? T_520_rd : T_407_rd;
  assign T_1846_rs1 = T_1655 ? T_520_rs1 : T_407_rs1;
  assign T_1846_rs2 = T_1655 ? T_520_rs2 : T_407_rs2;
  assign T_1846_rs3 = T_1655 ? T_520_rs3 : T_407_rs3;
  assign T_1852_bits = T_1651 ? T_1836_bits : T_1846_bits;
  assign T_1852_rd = T_1651 ? T_1836_rd : T_1846_rd;
  assign T_1852_rs1 = T_1651 ? T_1836_rs1 : T_1846_rs1;
  assign T_1852_rs2 = T_1651 ? T_1836_rs2 : T_1846_rs2;
  assign T_1852_rs3 = T_1651 ? T_1836_rs3 : T_1846_rs3;
  assign T_1858_bits = T_1647 ? T_1822_bits : T_1852_bits;
  assign T_1858_rd = T_1647 ? T_1822_rd : T_1852_rd;
  assign T_1858_rs1 = T_1647 ? T_1822_rs1 : T_1852_rs1;
  assign T_1858_rs2 = T_1647 ? T_1822_rs2 : T_1852_rs2;
  assign T_1858_rs3 = T_1647 ? T_1822_rs3 : T_1852_rs3;
  assign T_1876_bits = T_1655 ? T_374_bits : T_323_bits;
  assign T_1876_rd = T_1655 ? T_374_rd : T_323_rd;
  assign T_1876_rs1 = T_1655 ? T_374_rs1 : T_323_rs1;
  assign T_1876_rs2 = T_1655 ? T_374_rs2 : T_323_rs2;
  assign T_1876_rs3 = T_1655 ? T_374_rs3 : T_323_rs3;
  assign T_1886_bits = T_1655 ? T_272_bits : T_225_bits;
  assign T_1886_rd = T_1655 ? T_272_rd : T_225_rd;
  assign T_1886_rs1 = T_1655 ? T_272_rs1 : T_225_rs1;
  assign T_1886_rs2 = T_1655 ? T_272_rs2 : T_225_rs2;
  assign T_1886_rs3 = T_1655 ? T_272_rs3 : T_225_rs3;
  assign T_1892_bits = T_1651 ? T_1876_bits : T_1886_bits;
  assign T_1892_rd = T_1651 ? T_1876_rd : T_1886_rd;
  assign T_1892_rs1 = T_1651 ? T_1876_rs1 : T_1886_rs1;
  assign T_1892_rs2 = T_1651 ? T_1876_rs2 : T_1886_rs2;
  assign T_1892_rs3 = T_1651 ? T_1876_rs3 : T_1886_rs3;
  assign T_1906_bits = T_1655 ? T_174_bits : T_133_bits;
  assign T_1906_rd = T_1655 ? T_174_rd : T_133_rd;
  assign T_1906_rs1 = T_1655 ? T_174_rs1 : T_133_rs1;
  assign T_1906_rs2 = T_1655 ? T_174_rs2 : T_133_rs2;
  assign T_1906_rs3 = T_1655 ? T_174_rs3 : T_133_rs3;
  assign T_1916_bits = T_1655 ? T_92_bits : T_53_bits;
  assign T_1916_rd = T_1655 ? T_92_rd : T_53_rd;
  assign T_1916_rs1 = T_1655 ? T_92_rs1 : T_53_rs1;
  assign T_1916_rs2 = T_1655 ? T_92_rs2 : T_53_rs2;
  assign T_1916_rs3 = T_1655 ? T_92_rs3 : T_53_rs3;
  assign T_1922_bits = T_1651 ? T_1906_bits : T_1916_bits;
  assign T_1922_rd = T_1651 ? T_1906_rd : T_1916_rd;
  assign T_1922_rs1 = T_1651 ? T_1906_rs1 : T_1916_rs1;
  assign T_1922_rs2 = T_1651 ? T_1906_rs2 : T_1916_rs2;
  assign T_1922_rs3 = T_1651 ? T_1906_rs3 : T_1916_rs3;
  assign T_1928_bits = T_1647 ? T_1892_bits : T_1922_bits;
  assign T_1928_rd = T_1647 ? T_1892_rd : T_1922_rd;
  assign T_1928_rs1 = T_1647 ? T_1892_rs1 : T_1922_rs1;
  assign T_1928_rs2 = T_1647 ? T_1892_rs2 : T_1922_rs2;
  assign T_1928_rs3 = T_1647 ? T_1892_rs3 : T_1922_rs3;
  assign T_1934_bits = T_1643 ? T_1858_bits : T_1928_bits;
  assign T_1934_rd = T_1643 ? T_1858_rd : T_1928_rd;
  assign T_1934_rs1 = T_1643 ? T_1858_rs1 : T_1928_rs1;
  assign T_1934_rs2 = T_1643 ? T_1858_rs2 : T_1928_rs2;
  assign T_1934_rs3 = T_1643 ? T_1858_rs3 : T_1928_rs3;
  assign T_1940_bits = T_1639 ? T_1784_bits : T_1934_bits;
  assign T_1940_rd = T_1639 ? T_1784_rd : T_1934_rd;
  assign T_1940_rs1 = T_1639 ? T_1784_rs1 : T_1934_rs1;
  assign T_1940_rs2 = T_1639 ? T_1784_rs2 : T_1934_rs2;
  assign T_1940_rs3 = T_1639 ? T_1784_rs3 : T_1934_rs3;
endmodule