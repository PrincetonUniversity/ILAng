/* PREHEADER */
module fun_gb_fun (
    input [647:0] arg1,
    output [7:0] result
);
//TODO: Add the specific function HERE.
endmodule

/* END OF PREHEADER */
module SPEC_A(
arg_0_TREADY,
arg_1_TDATA,
arg_1_TVALID,
RAM_w,
RAM_x,
RAM_y,
arg_0_TDATA,
arg_0_TVALID,
arg_1_TREADY,
cur_pix,
gbit,
pre_pix,
proc_in,
st_ready,
stencil_0,
stencil_1,
stencil_2,
stencil_3,
stencil_4,
stencil_5,
stencil_6,
stencil_7,
stencil_8,
clk,rst,
step
);
input            arg_0_TREADY;
input      [7:0] arg_1_TDATA;
input            arg_1_TVALID;
input clk;
input rst;
input step;
output      [2:0] RAM_w;
output      [8:0] RAM_x;
output      [9:0] RAM_y;
output      [7:0] arg_0_TDATA;
output            arg_0_TVALID;
output            arg_1_TREADY;
output      [7:0] cur_pix;
output      [3:0] gbit;
output      [7:0] pre_pix;
output    [647:0] proc_in;
output            st_ready;
output     [71:0] stencil_0;
output     [71:0] stencil_1;
output     [71:0] stencil_2;
output     [71:0] stencil_3;
output     [71:0] stencil_4;
output     [71:0] stencil_5;
output     [71:0] stencil_6;
output     [71:0] stencil_7;
output     [71:0] stencil_8;
reg      [2:0] RAM_w;
reg      [8:0] RAM_x;
reg      [9:0] RAM_y;
reg      [7:0] arg_0_TDATA;
reg            arg_0_TVALID;
reg            arg_1_TREADY;
reg      [7:0] cur_pix;
reg      [3:0] gbit;
reg      [7:0] pre_pix;
reg    [647:0] proc_in;
reg            st_ready;
reg     [71:0] stencil_0;
reg     [71:0] stencil_1;
reg     [71:0] stencil_2;
reg     [71:0] stencil_3;
reg     [71:0] stencil_4;
reg     [71:0] stencil_5;
reg     [71:0] stencil_6;
reg     [71:0] stencil_7;
reg     [71:0] stencil_8;
wire            arg_0_TREADY;
wire      [7:0] arg_1_TDATA;
wire            arg_1_TVALID;
wire            n0;
wire            n1;
wire            n2;
wire            n3;
wire            n4;
wire            n5;
wire            n6;
wire            n7;
wire            n8;
wire      [2:0] n9;
wire      [2:0] n10;
wire      [2:0] n11;
wire            n12;
wire            n13;
wire            n14;
wire            n15;
wire            n16;
wire            n17;
wire      [2:0] n18;
wire      [2:0] n19;
wire      [2:0] n20;
wire            n21;
wire            n22;
wire            n23;
wire      [8:0] n24;
wire      [8:0] n25;
wire      [8:0] n26;
wire      [8:0] n27;
wire      [8:0] n28;
wire      [8:0] n29;
wire            n30;
wire      [9:0] n31;
wire      [9:0] n32;
wire      [9:0] n33;
wire      [9:0] n34;
wire      [9:0] n35;
wire      [9:0] n36;
wire            n37;
wire            n38;
wire            n39;
wire            n40;
wire            n41;
wire            n42;
wire            n43;
wire            n44;
wire      [7:0] n45;
wire      [7:0] n46;
wire      [7:0] n47;
wire      [7:0] n48;
wire      [7:0] n49;
wire      [7:0] n50;
wire      [7:0] n51;
wire      [7:0] n52;
wire      [7:0] n53;
wire     [15:0] n54;
wire     [23:0] n55;
wire     [31:0] n56;
wire     [39:0] n57;
wire     [47:0] n58;
wire     [55:0] n59;
wire     [63:0] n60;
wire     [71:0] n61;
wire      [7:0] n62;
wire      [7:0] n63;
wire      [7:0] n64;
wire      [7:0] n65;
wire      [7:0] n66;
wire      [7:0] n67;
wire      [7:0] n68;
wire      [7:0] n69;
wire      [7:0] n70;
wire     [15:0] n71;
wire     [23:0] n72;
wire     [31:0] n73;
wire     [39:0] n74;
wire     [47:0] n75;
wire     [55:0] n76;
wire     [63:0] n77;
wire     [71:0] n78;
wire      [7:0] n79;
wire      [7:0] n80;
wire      [7:0] n81;
wire      [7:0] n82;
wire      [7:0] n83;
wire      [7:0] n84;
wire      [7:0] n85;
wire      [7:0] n86;
wire      [7:0] n87;
wire     [15:0] n88;
wire     [23:0] n89;
wire     [31:0] n90;
wire     [39:0] n91;
wire     [47:0] n92;
wire     [55:0] n93;
wire     [63:0] n94;
wire     [71:0] n95;
wire      [7:0] n96;
wire      [7:0] n97;
wire      [7:0] n98;
wire      [7:0] n99;
wire      [7:0] n100;
wire      [7:0] n101;
wire      [7:0] n102;
wire      [7:0] n103;
wire      [7:0] n104;
wire     [15:0] n105;
wire     [23:0] n106;
wire     [31:0] n107;
wire     [39:0] n108;
wire     [47:0] n109;
wire     [55:0] n110;
wire     [63:0] n111;
wire     [71:0] n112;
wire      [7:0] n113;
wire      [7:0] n114;
wire      [7:0] n115;
wire      [7:0] n116;
wire      [7:0] n117;
wire      [7:0] n118;
wire      [7:0] n119;
wire      [7:0] n120;
wire      [7:0] n121;
wire     [15:0] n122;
wire     [23:0] n123;
wire     [31:0] n124;
wire     [39:0] n125;
wire     [47:0] n126;
wire     [55:0] n127;
wire     [63:0] n128;
wire     [71:0] n129;
wire      [7:0] n130;
wire      [7:0] n131;
wire      [7:0] n132;
wire      [7:0] n133;
wire      [7:0] n134;
wire      [7:0] n135;
wire      [7:0] n136;
wire      [7:0] n137;
wire      [7:0] n138;
wire     [15:0] n139;
wire     [23:0] n140;
wire     [31:0] n141;
wire     [39:0] n142;
wire     [47:0] n143;
wire     [55:0] n144;
wire     [63:0] n145;
wire     [71:0] n146;
wire      [7:0] n147;
wire      [7:0] n148;
wire      [7:0] n149;
wire      [7:0] n150;
wire      [7:0] n151;
wire      [7:0] n152;
wire      [7:0] n153;
wire      [7:0] n154;
wire      [7:0] n155;
wire     [15:0] n156;
wire     [23:0] n157;
wire     [31:0] n158;
wire     [39:0] n159;
wire     [47:0] n160;
wire     [55:0] n161;
wire     [63:0] n162;
wire     [71:0] n163;
wire      [7:0] n164;
wire      [7:0] n165;
wire      [7:0] n166;
wire      [7:0] n167;
wire      [7:0] n168;
wire      [7:0] n169;
wire      [7:0] n170;
wire      [7:0] n171;
wire      [7:0] n172;
wire     [15:0] n173;
wire     [23:0] n174;
wire     [31:0] n175;
wire     [39:0] n176;
wire     [47:0] n177;
wire     [55:0] n178;
wire     [63:0] n179;
wire     [71:0] n180;
wire      [7:0] n181;
wire      [7:0] n182;
wire      [7:0] n183;
wire      [7:0] n184;
wire      [7:0] n185;
wire      [7:0] n186;
wire      [7:0] n187;
wire      [7:0] n188;
wire      [7:0] n189;
wire     [15:0] n190;
wire     [23:0] n191;
wire     [31:0] n192;
wire     [39:0] n193;
wire     [47:0] n194;
wire     [55:0] n195;
wire     [63:0] n196;
wire     [71:0] n197;
wire    [143:0] n198;
wire    [215:0] n199;
wire    [287:0] n200;
wire    [359:0] n201;
wire    [431:0] n202;
wire    [503:0] n203;
wire    [575:0] n204;
wire    [647:0] n205;
wire    [647:0] n206;
wire    [647:0] n207;
wire      [7:0] n208;
wire      [7:0] n210;
wire      [7:0] n211;
wire      [7:0] n212;
wire      [7:0] n213;
wire      [7:0] n214;
wire            n215;
wire            n216;
wire            n217;
wire            n218;
wire            n219;
wire            n220;
wire      [8:0] n221;
wire            n222;
wire      [9:0] n223;
wire            n224;
wire            n225;
wire            n226;
wire            n227;
wire            n228;
wire            n229;
wire            n230;
wire            n231;
wire            n232;
wire      [7:0] n233;
wire      [7:0] n234;
wire      [7:0] n235;
wire      [7:0] n236;
wire      [7:0] n237;
wire    [647:0] n238;
wire    [647:0] n239;
wire            n240;
wire            n241;
wire     [71:0] n242;
wire     [71:0] n243;
wire     [71:0] n244;
wire     [71:0] n245;
wire     [71:0] n246;
wire     [71:0] n247;
wire     [71:0] n248;
wire     [71:0] n249;
wire     [71:0] n250;
wire     [71:0] n251;
wire     [71:0] n252;
wire     [71:0] n253;
wire     [71:0] n254;
wire     [71:0] n255;
wire     [71:0] n256;
wire     [71:0] n257;
wire     [71:0] n258;
wire     [71:0] n259;
wire     [71:0] n260;
wire     [71:0] n261;
wire     [71:0] n262;
wire     [71:0] n263;
wire     [71:0] n264;
wire     [71:0] n265;
wire     [71:0] n266;
wire     [71:0] n267;
wire     [71:0] n268;
wire     [71:0] n269;
wire     [71:0] n270;
wire     [71:0] n271;
wire     [71:0] n272;
wire     [71:0] n273;
wire            n274;
wire      [8:0] n275;
wire      [7:0] n276;
wire            n277;
wire      [7:0] n278;
wire            n279;
wire      [7:0] n280;
wire            n281;
wire      [7:0] n282;
wire            n283;
wire      [7:0] n284;
wire            n285;
wire      [7:0] n286;
wire            n287;
wire      [7:0] n288;
wire      [7:0] n289;
wire      [7:0] n290;
wire      [7:0] n291;
wire      [7:0] n292;
wire      [7:0] n293;
wire      [7:0] n294;
wire      [7:0] n295;
wire      [7:0] n296;
wire      [7:0] n297;
wire      [7:0] n298;
wire      [7:0] n299;
wire      [7:0] n300;
wire      [7:0] n301;
wire      [7:0] n302;
wire      [7:0] n303;
wire      [7:0] n304;
wire      [7:0] n305;
wire      [7:0] n306;
wire      [7:0] n307;
wire      [7:0] n308;
wire      [7:0] n309;
wire      [7:0] n310;
wire      [7:0] n311;
wire      [7:0] n312;
wire      [7:0] n313;
wire      [7:0] n314;
wire      [7:0] n315;
wire      [7:0] n316;
wire      [7:0] n317;
wire      [7:0] n318;
wire      [7:0] n319;
wire      [7:0] n320;
wire      [7:0] n321;
wire      [7:0] n322;
wire      [7:0] n323;
wire      [7:0] n324;
wire      [7:0] n325;
wire      [7:0] n326;
wire      [7:0] n327;
wire      [7:0] n328;
wire      [7:0] n329;
wire      [7:0] n330;
wire      [7:0] n331;
wire      [7:0] n332;
wire      [7:0] n333;
wire      [7:0] n334;
wire      [7:0] n335;
wire      [7:0] n336;
wire      [7:0] n337;
wire      [7:0] n338;
wire      [7:0] n339;
wire      [7:0] n340;
wire      [7:0] n341;
wire      [7:0] n342;
wire      [7:0] n343;
wire      [7:0] n344;
wire      [7:0] n345;
wire     [15:0] n346;
wire     [23:0] n347;
wire     [31:0] n348;
wire     [39:0] n349;
wire     [47:0] n350;
wire     [55:0] n351;
wire     [63:0] n352;
wire     [71:0] n353;
wire     [71:0] n354;
wire     [71:0] n355;
wire     [71:0] n356;
wire     [71:0] n357;
wire      [8:0] RAM_0_addr0;
wire      [7:0] RAM_0_data0;
wire            RAM_0_wen0;
wire            n358;
wire            n359;
wire            n360;
wire            n361;
wire            n362;
wire            n363;
wire            n364;
wire            n365;
wire            n366;
wire            n367;
wire            n368;
wire            n369;
wire            n370;
wire            n371;
wire            n372;
wire      [8:0] RAM_1_addr0;
wire      [7:0] RAM_1_data0;
wire            RAM_1_wen0;
wire            n373;
wire            n374;
wire            n375;
wire      [8:0] RAM_2_addr0;
wire      [7:0] RAM_2_data0;
wire            RAM_2_wen0;
wire            n376;
wire            n377;
wire            n378;
wire      [8:0] RAM_3_addr0;
wire      [7:0] RAM_3_data0;
wire            RAM_3_wen0;
wire            n379;
wire            n380;
wire            n381;
wire      [8:0] RAM_4_addr0;
wire      [7:0] RAM_4_data0;
wire            RAM_4_wen0;
wire            n382;
wire            n383;
wire            n384;
wire      [8:0] RAM_5_addr0;
wire      [7:0] RAM_5_data0;
wire            RAM_5_wen0;
wire            n385;
wire            n386;
wire            n387;
wire      [8:0] RAM_6_addr0;
wire      [7:0] RAM_6_data0;
wire            RAM_6_wen0;
wire            n388;
wire            n389;
wire            n390;
wire      [8:0] RAM_7_addr0;
wire      [7:0] RAM_7_data0;
wire            RAM_7_wen0;
wire            n391;
wire            n392;
wire            n393;
reg      [7:0] RAM_0[487:0];
reg      [7:0] RAM_1[487:0];
reg      [7:0] RAM_2[487:0];
reg      [7:0] RAM_3[487:0];
reg      [7:0] RAM_4[487:0];
reg      [7:0] RAM_5[487:0];
reg      [7:0] RAM_6[487:0];
reg      [7:0] RAM_7[487:0];
wire clk;
wire rst;
wire step;
assign n0 =  ( arg_1_TREADY ) == ( 1'd0 )  ;
assign n1 =  ( arg_0_TREADY ) == ( 1'd0 )  ;
assign n2 =  ( n0 ) & ( n1 )  ;
assign n3 =  ( st_ready ) == ( 1'd0 )  ;
assign n4 =  ( n2 ) & ( n3 )  ;
assign n5 =  ( st_ready ) == ( 1'd1 )  ;
assign n6 =  ( n2 ) & ( n5 )  ;
assign n7 =  ( RAM_x ) == ( 9'd488 )  ;
assign n8 =  ( RAM_w ) == ( 3'd7 )  ;
assign n9 =  ( RAM_w ) + ( 3'd1 )  ;
assign n10 =  ( n8 ) ? ( 3'd0 ) : ( n9 ) ;
assign n11 =  ( n7 ) ? ( n10 ) : ( RAM_w ) ;
assign n12 =  ( arg_1_TVALID ) == ( 1'd1 )  ;
assign n13 =  ( arg_1_TREADY ) == ( 1'd1 )  ;
assign n14 =  ( n12 ) & ( n13 )  ;
assign n15 =  ( arg_0_TVALID ) == ( 1'd0 )  ;
assign n16 =  ( n14 ) & ( n15 )  ;
assign n17 =  ( n16 ) & ( n1 )  ;
assign n18 =  ( n17 ) ? ( RAM_w ) : ( RAM_w ) ;
assign n19 =  ( n6 ) ? ( n11 ) : ( n18 ) ;
assign n20 =  ( n4 ) ? ( RAM_w ) : ( n19 ) ;
assign n21 =  ( RAM_x ) == ( 9'd0 )  ;
assign n22 =  ( RAM_y ) == ( 10'd0 )  ;
assign n23 =  ( n21 ) & ( n22 )  ;
assign n24 =  ( RAM_x ) + ( 9'd1 )  ;
assign n25 =  ( n7 ) ? ( 9'd1 ) : ( n24 ) ;
assign n26 =  ( n23 ) ? ( 9'd1 ) : ( n25 ) ;
assign n27 =  ( n17 ) ? ( RAM_x ) : ( RAM_x ) ;
assign n28 =  ( n6 ) ? ( n26 ) : ( n27 ) ;
assign n29 =  ( n4 ) ? ( RAM_x ) : ( n28 ) ;
assign n30 =  ( RAM_y ) == ( 10'd648 )  ;
assign n31 =  ( RAM_y ) + ( 10'd1 )  ;
assign n32 =  ( n30 ) ? ( 10'd0 ) : ( n31 ) ;
assign n33 =  ( n7 ) ? ( n32 ) : ( RAM_y ) ;
assign n34 =  ( n17 ) ? ( RAM_y ) : ( RAM_y ) ;
assign n35 =  ( n6 ) ? ( n33 ) : ( n34 ) ;
assign n36 =  ( n4 ) ? ( RAM_y ) : ( n35 ) ;
assign n37 =  ( RAM_x ) == ( 9'd1 )  ;
assign n38 =  ( n37 ) & ( n30 )  ;
assign n39 =  ( RAM_x ) > ( 9'd8 )  ;
assign n40 =  ( RAM_y ) >= ( 10'd8 )  ;
assign n41 =  ( n39 ) & ( n40 )  ;
assign n42 =  ( RAM_y ) > ( 10'd8 )  ;
assign n43 =  ( n37 ) & ( n42 )  ;
assign n44 =  ( n41 ) | ( n43 )  ;
assign n45 = stencil_8[71:64] ;
assign n46 = stencil_7[71:64] ;
assign n47 = stencil_6[71:64] ;
assign n48 = stencil_5[71:64] ;
assign n49 = stencil_4[71:64] ;
assign n50 = stencil_3[71:64] ;
assign n51 = stencil_2[71:64] ;
assign n52 = stencil_1[71:64] ;
assign n53 = stencil_0[71:64] ;
assign n54 =  { ( n52 ) , ( n53 ) }  ;
assign n55 =  { ( n51 ) , ( n54 ) }  ;
assign n56 =  { ( n50 ) , ( n55 ) }  ;
assign n57 =  { ( n49 ) , ( n56 ) }  ;
assign n58 =  { ( n48 ) , ( n57 ) }  ;
assign n59 =  { ( n47 ) , ( n58 ) }  ;
assign n60 =  { ( n46 ) , ( n59 ) }  ;
assign n61 =  { ( n45 ) , ( n60 ) }  ;
assign n62 = stencil_8[63:56] ;
assign n63 = stencil_7[63:56] ;
assign n64 = stencil_6[63:56] ;
assign n65 = stencil_5[63:56] ;
assign n66 = stencil_4[63:56] ;
assign n67 = stencil_3[63:56] ;
assign n68 = stencil_2[63:56] ;
assign n69 = stencil_1[63:56] ;
assign n70 = stencil_0[63:56] ;
assign n71 =  { ( n69 ) , ( n70 ) }  ;
assign n72 =  { ( n68 ) , ( n71 ) }  ;
assign n73 =  { ( n67 ) , ( n72 ) }  ;
assign n74 =  { ( n66 ) , ( n73 ) }  ;
assign n75 =  { ( n65 ) , ( n74 ) }  ;
assign n76 =  { ( n64 ) , ( n75 ) }  ;
assign n77 =  { ( n63 ) , ( n76 ) }  ;
assign n78 =  { ( n62 ) , ( n77 ) }  ;
assign n79 = stencil_8[55:48] ;
assign n80 = stencil_7[55:48] ;
assign n81 = stencil_6[55:48] ;
assign n82 = stencil_5[55:48] ;
assign n83 = stencil_4[55:48] ;
assign n84 = stencil_3[55:48] ;
assign n85 = stencil_2[55:48] ;
assign n86 = stencil_1[55:48] ;
assign n87 = stencil_0[55:48] ;
assign n88 =  { ( n86 ) , ( n87 ) }  ;
assign n89 =  { ( n85 ) , ( n88 ) }  ;
assign n90 =  { ( n84 ) , ( n89 ) }  ;
assign n91 =  { ( n83 ) , ( n90 ) }  ;
assign n92 =  { ( n82 ) , ( n91 ) }  ;
assign n93 =  { ( n81 ) , ( n92 ) }  ;
assign n94 =  { ( n80 ) , ( n93 ) }  ;
assign n95 =  { ( n79 ) , ( n94 ) }  ;
assign n96 = stencil_8[47:40] ;
assign n97 = stencil_7[47:40] ;
assign n98 = stencil_6[47:40] ;
assign n99 = stencil_5[47:40] ;
assign n100 = stencil_4[47:40] ;
assign n101 = stencil_3[47:40] ;
assign n102 = stencil_2[47:40] ;
assign n103 = stencil_1[47:40] ;
assign n104 = stencil_0[47:40] ;
assign n105 =  { ( n103 ) , ( n104 ) }  ;
assign n106 =  { ( n102 ) , ( n105 ) }  ;
assign n107 =  { ( n101 ) , ( n106 ) }  ;
assign n108 =  { ( n100 ) , ( n107 ) }  ;
assign n109 =  { ( n99 ) , ( n108 ) }  ;
assign n110 =  { ( n98 ) , ( n109 ) }  ;
assign n111 =  { ( n97 ) , ( n110 ) }  ;
assign n112 =  { ( n96 ) , ( n111 ) }  ;
assign n113 = stencil_8[39:32] ;
assign n114 = stencil_7[39:32] ;
assign n115 = stencil_6[39:32] ;
assign n116 = stencil_5[39:32] ;
assign n117 = stencil_4[39:32] ;
assign n118 = stencil_3[39:32] ;
assign n119 = stencil_2[39:32] ;
assign n120 = stencil_1[39:32] ;
assign n121 = stencil_0[39:32] ;
assign n122 =  { ( n120 ) , ( n121 ) }  ;
assign n123 =  { ( n119 ) , ( n122 ) }  ;
assign n124 =  { ( n118 ) , ( n123 ) }  ;
assign n125 =  { ( n117 ) , ( n124 ) }  ;
assign n126 =  { ( n116 ) , ( n125 ) }  ;
assign n127 =  { ( n115 ) , ( n126 ) }  ;
assign n128 =  { ( n114 ) , ( n127 ) }  ;
assign n129 =  { ( n113 ) , ( n128 ) }  ;
assign n130 = stencil_8[31:24] ;
assign n131 = stencil_7[31:24] ;
assign n132 = stencil_6[31:24] ;
assign n133 = stencil_5[31:24] ;
assign n134 = stencil_4[31:24] ;
assign n135 = stencil_3[31:24] ;
assign n136 = stencil_2[31:24] ;
assign n137 = stencil_1[31:24] ;
assign n138 = stencil_0[31:24] ;
assign n139 =  { ( n137 ) , ( n138 ) }  ;
assign n140 =  { ( n136 ) , ( n139 ) }  ;
assign n141 =  { ( n135 ) , ( n140 ) }  ;
assign n142 =  { ( n134 ) , ( n141 ) }  ;
assign n143 =  { ( n133 ) , ( n142 ) }  ;
assign n144 =  { ( n132 ) , ( n143 ) }  ;
assign n145 =  { ( n131 ) , ( n144 ) }  ;
assign n146 =  { ( n130 ) , ( n145 ) }  ;
assign n147 = stencil_8[23:16] ;
assign n148 = stencil_7[23:16] ;
assign n149 = stencil_6[23:16] ;
assign n150 = stencil_5[23:16] ;
assign n151 = stencil_4[23:16] ;
assign n152 = stencil_3[23:16] ;
assign n153 = stencil_2[23:16] ;
assign n154 = stencil_1[23:16] ;
assign n155 = stencil_0[23:16] ;
assign n156 =  { ( n154 ) , ( n155 ) }  ;
assign n157 =  { ( n153 ) , ( n156 ) }  ;
assign n158 =  { ( n152 ) , ( n157 ) }  ;
assign n159 =  { ( n151 ) , ( n158 ) }  ;
assign n160 =  { ( n150 ) , ( n159 ) }  ;
assign n161 =  { ( n149 ) , ( n160 ) }  ;
assign n162 =  { ( n148 ) , ( n161 ) }  ;
assign n163 =  { ( n147 ) , ( n162 ) }  ;
assign n164 = stencil_8[15:8] ;
assign n165 = stencil_7[15:8] ;
assign n166 = stencil_6[15:8] ;
assign n167 = stencil_5[15:8] ;
assign n168 = stencil_4[15:8] ;
assign n169 = stencil_3[15:8] ;
assign n170 = stencil_2[15:8] ;
assign n171 = stencil_1[15:8] ;
assign n172 = stencil_0[15:8] ;
assign n173 =  { ( n171 ) , ( n172 ) }  ;
assign n174 =  { ( n170 ) , ( n173 ) }  ;
assign n175 =  { ( n169 ) , ( n174 ) }  ;
assign n176 =  { ( n168 ) , ( n175 ) }  ;
assign n177 =  { ( n167 ) , ( n176 ) }  ;
assign n178 =  { ( n166 ) , ( n177 ) }  ;
assign n179 =  { ( n165 ) , ( n178 ) }  ;
assign n180 =  { ( n164 ) , ( n179 ) }  ;
assign n181 = stencil_8[7:0] ;
assign n182 = stencil_7[7:0] ;
assign n183 = stencil_6[7:0] ;
assign n184 = stencil_5[7:0] ;
assign n185 = stencil_4[7:0] ;
assign n186 = stencil_3[7:0] ;
assign n187 = stencil_2[7:0] ;
assign n188 = stencil_1[7:0] ;
assign n189 = stencil_0[7:0] ;
assign n190 =  { ( n188 ) , ( n189 ) }  ;
assign n191 =  { ( n187 ) , ( n190 ) }  ;
assign n192 =  { ( n186 ) , ( n191 ) }  ;
assign n193 =  { ( n185 ) , ( n192 ) }  ;
assign n194 =  { ( n184 ) , ( n193 ) }  ;
assign n195 =  { ( n183 ) , ( n194 ) }  ;
assign n196 =  { ( n182 ) , ( n195 ) }  ;
assign n197 =  { ( n181 ) , ( n196 ) }  ;
assign n198 =  { ( n180 ) , ( n197 ) }  ;
assign n199 =  { ( n163 ) , ( n198 ) }  ;
assign n200 =  { ( n146 ) , ( n199 ) }  ;
assign n201 =  { ( n129 ) , ( n200 ) }  ;
assign n202 =  { ( n112 ) , ( n201 ) }  ;
assign n203 =  { ( n95 ) , ( n202 ) }  ;
assign n204 =  { ( n78 ) , ( n203 ) }  ;
assign n205 =  { ( n61 ) , ( n204 ) }  ;
assign n206 =  ( n44 ) ? ( n205 ) : ( proc_in ) ;
assign n207 =  ( n38 ) ? ( proc_in ) : ( n206 ) ;
fun_gb_fun  applyFunc_n209(
    .arg1( n207 ),
    .result( n208 )
);
assign n210 = n208 ;
assign n211 =  ( n38 ) ? ( arg_0_TDATA ) : ( n210 ) ;
assign n212 =  ( n17 ) ? ( arg_0_TDATA ) : ( arg_0_TDATA ) ;
assign n213 =  ( n6 ) ? ( arg_0_TDATA ) : ( n212 ) ;
assign n214 =  ( n4 ) ? ( n211 ) : ( n213 ) ;
assign n215 =  ( n44 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n216 =  ( n38 ) ? ( arg_0_TVALID ) : ( n215 ) ;
assign n217 =  ( n23 ) ? ( 1'd0 ) : ( arg_0_TVALID ) ;
assign n218 =  ( n17 ) ? ( 1'd0 ) : ( arg_0_TVALID ) ;
assign n219 =  ( n6 ) ? ( n217 ) : ( n218 ) ;
assign n220 =  ( n4 ) ? ( n216 ) : ( n219 ) ;
assign n221 =  ( 9'd488 ) - ( 9'd1 )  ;
assign n222 =  ( RAM_x ) == ( n221 )  ;
assign n223 =  ( 10'd648 ) - ( 10'd1 )  ;
assign n224 =  ( RAM_y ) == ( n223 )  ;
assign n225 =  ( n222 ) & ( n224 )  ;
assign n226 =  ( n225 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n227 =  ( RAM_y ) < ( 10'd8 )  ;
assign n228 =  ( n227 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n229 =  ( n23 ) ? ( 1'd1 ) : ( n228 ) ;
assign n230 =  ( n17 ) ? ( 1'd0 ) : ( arg_1_TREADY ) ;
assign n231 =  ( n6 ) ? ( n229 ) : ( n230 ) ;
assign n232 =  ( n4 ) ? ( n226 ) : ( n231 ) ;
assign n233 =  ( n17 ) ? ( arg_1_TDATA ) : ( cur_pix ) ;
assign n234 =  ( n6 ) ? ( cur_pix ) : ( n233 ) ;
assign n235 =  ( n4 ) ? ( cur_pix ) : ( n234 ) ;
assign n236 =  ( n6 ) ? ( cur_pix ) : ( pre_pix ) ;
assign n237 =  ( n4 ) ? ( pre_pix ) : ( n236 ) ;
assign n238 =  ( n6 ) ? ( proc_in ) : ( proc_in ) ;
assign n239 =  ( n4 ) ? ( n207 ) : ( n238 ) ;
assign n240 =  ( n6 ) ? ( n229 ) : ( st_ready ) ;
assign n241 =  ( n4 ) ? ( 1'd1 ) : ( n240 ) ;
assign n242 =  ( n227 ) ? ( stencil_0 ) : ( stencil_1 ) ;
assign n243 =  ( n17 ) ? ( stencil_0 ) : ( stencil_0 ) ;
assign n244 =  ( n6 ) ? ( stencil_0 ) : ( n243 ) ;
assign n245 =  ( n4 ) ? ( n242 ) : ( n244 ) ;
assign n246 =  ( n227 ) ? ( stencil_1 ) : ( stencil_2 ) ;
assign n247 =  ( n17 ) ? ( stencil_1 ) : ( stencil_1 ) ;
assign n248 =  ( n6 ) ? ( stencil_1 ) : ( n247 ) ;
assign n249 =  ( n4 ) ? ( n246 ) : ( n248 ) ;
assign n250 =  ( n227 ) ? ( stencil_2 ) : ( stencil_3 ) ;
assign n251 =  ( n17 ) ? ( stencil_2 ) : ( stencil_2 ) ;
assign n252 =  ( n6 ) ? ( stencil_2 ) : ( n251 ) ;
assign n253 =  ( n4 ) ? ( n250 ) : ( n252 ) ;
assign n254 =  ( n227 ) ? ( stencil_3 ) : ( stencil_4 ) ;
assign n255 =  ( n17 ) ? ( stencil_3 ) : ( stencil_3 ) ;
assign n256 =  ( n6 ) ? ( stencil_3 ) : ( n255 ) ;
assign n257 =  ( n4 ) ? ( n254 ) : ( n256 ) ;
assign n258 =  ( n227 ) ? ( stencil_4 ) : ( stencil_5 ) ;
assign n259 =  ( n17 ) ? ( stencil_4 ) : ( stencil_4 ) ;
assign n260 =  ( n6 ) ? ( stencil_4 ) : ( n259 ) ;
assign n261 =  ( n4 ) ? ( n258 ) : ( n260 ) ;
assign n262 =  ( n227 ) ? ( stencil_5 ) : ( stencil_6 ) ;
assign n263 =  ( n17 ) ? ( stencil_5 ) : ( stencil_5 ) ;
assign n264 =  ( n6 ) ? ( stencil_5 ) : ( n263 ) ;
assign n265 =  ( n4 ) ? ( n262 ) : ( n264 ) ;
assign n266 =  ( n227 ) ? ( stencil_6 ) : ( stencil_7 ) ;
assign n267 =  ( n17 ) ? ( stencil_6 ) : ( stencil_6 ) ;
assign n268 =  ( n6 ) ? ( stencil_6 ) : ( n267 ) ;
assign n269 =  ( n4 ) ? ( n266 ) : ( n268 ) ;
assign n270 =  ( n227 ) ? ( stencil_7 ) : ( stencil_8 ) ;
assign n271 =  ( n17 ) ? ( stencil_7 ) : ( stencil_7 ) ;
assign n272 =  ( n6 ) ? ( stencil_7 ) : ( n271 ) ;
assign n273 =  ( n4 ) ? ( n270 ) : ( n272 ) ;
assign n274 =  ( RAM_w ) == ( 3'd0 )  ;
assign n275 =  ( RAM_x ) - ( 9'd1 )  ;
assign n276 =  (  RAM_7 [ n275 ] )  ;
assign n277 =  ( RAM_w ) == ( 3'd1 )  ;
assign n278 =  (  RAM_0 [ n275 ] )  ;
assign n279 =  ( RAM_w ) == ( 3'd2 )  ;
assign n280 =  (  RAM_1 [ n275 ] )  ;
assign n281 =  ( RAM_w ) == ( 3'd3 )  ;
assign n282 =  (  RAM_2 [ n275 ] )  ;
assign n283 =  ( RAM_w ) == ( 3'd4 )  ;
assign n284 =  (  RAM_3 [ n275 ] )  ;
assign n285 =  ( RAM_w ) == ( 3'd5 )  ;
assign n286 =  (  RAM_4 [ n275 ] )  ;
assign n287 =  ( RAM_w ) == ( 3'd6 )  ;
assign n288 =  (  RAM_5 [ n275 ] )  ;
assign n289 =  (  RAM_6 [ n275 ] )  ;
assign n290 =  ( n287 ) ? ( n288 ) : ( n289 ) ;
assign n291 =  ( n285 ) ? ( n286 ) : ( n290 ) ;
assign n292 =  ( n283 ) ? ( n284 ) : ( n291 ) ;
assign n293 =  ( n281 ) ? ( n282 ) : ( n292 ) ;
assign n294 =  ( n279 ) ? ( n280 ) : ( n293 ) ;
assign n295 =  ( n277 ) ? ( n278 ) : ( n294 ) ;
assign n296 =  ( n274 ) ? ( n276 ) : ( n295 ) ;
assign n297 =  ( n287 ) ? ( n286 ) : ( n288 ) ;
assign n298 =  ( n285 ) ? ( n284 ) : ( n297 ) ;
assign n299 =  ( n283 ) ? ( n282 ) : ( n298 ) ;
assign n300 =  ( n281 ) ? ( n280 ) : ( n299 ) ;
assign n301 =  ( n279 ) ? ( n278 ) : ( n300 ) ;
assign n302 =  ( n277 ) ? ( n276 ) : ( n301 ) ;
assign n303 =  ( n274 ) ? ( n289 ) : ( n302 ) ;
assign n304 =  ( n287 ) ? ( n284 ) : ( n286 ) ;
assign n305 =  ( n285 ) ? ( n282 ) : ( n304 ) ;
assign n306 =  ( n283 ) ? ( n280 ) : ( n305 ) ;
assign n307 =  ( n281 ) ? ( n278 ) : ( n306 ) ;
assign n308 =  ( n279 ) ? ( n276 ) : ( n307 ) ;
assign n309 =  ( n277 ) ? ( n289 ) : ( n308 ) ;
assign n310 =  ( n274 ) ? ( n288 ) : ( n309 ) ;
assign n311 =  ( n287 ) ? ( n282 ) : ( n284 ) ;
assign n312 =  ( n285 ) ? ( n280 ) : ( n311 ) ;
assign n313 =  ( n283 ) ? ( n278 ) : ( n312 ) ;
assign n314 =  ( n281 ) ? ( n276 ) : ( n313 ) ;
assign n315 =  ( n279 ) ? ( n289 ) : ( n314 ) ;
assign n316 =  ( n277 ) ? ( n288 ) : ( n315 ) ;
assign n317 =  ( n274 ) ? ( n286 ) : ( n316 ) ;
assign n318 =  ( n287 ) ? ( n280 ) : ( n282 ) ;
assign n319 =  ( n285 ) ? ( n278 ) : ( n318 ) ;
assign n320 =  ( n283 ) ? ( n276 ) : ( n319 ) ;
assign n321 =  ( n281 ) ? ( n289 ) : ( n320 ) ;
assign n322 =  ( n279 ) ? ( n288 ) : ( n321 ) ;
assign n323 =  ( n277 ) ? ( n286 ) : ( n322 ) ;
assign n324 =  ( n274 ) ? ( n284 ) : ( n323 ) ;
assign n325 =  ( n287 ) ? ( n278 ) : ( n280 ) ;
assign n326 =  ( n285 ) ? ( n276 ) : ( n325 ) ;
assign n327 =  ( n283 ) ? ( n289 ) : ( n326 ) ;
assign n328 =  ( n281 ) ? ( n288 ) : ( n327 ) ;
assign n329 =  ( n279 ) ? ( n286 ) : ( n328 ) ;
assign n330 =  ( n277 ) ? ( n284 ) : ( n329 ) ;
assign n331 =  ( n274 ) ? ( n282 ) : ( n330 ) ;
assign n332 =  ( n287 ) ? ( n276 ) : ( n278 ) ;
assign n333 =  ( n285 ) ? ( n289 ) : ( n332 ) ;
assign n334 =  ( n283 ) ? ( n288 ) : ( n333 ) ;
assign n335 =  ( n281 ) ? ( n286 ) : ( n334 ) ;
assign n336 =  ( n279 ) ? ( n284 ) : ( n335 ) ;
assign n337 =  ( n277 ) ? ( n282 ) : ( n336 ) ;
assign n338 =  ( n274 ) ? ( n280 ) : ( n337 ) ;
assign n339 =  ( n287 ) ? ( n289 ) : ( n276 ) ;
assign n340 =  ( n285 ) ? ( n288 ) : ( n339 ) ;
assign n341 =  ( n283 ) ? ( n286 ) : ( n340 ) ;
assign n342 =  ( n281 ) ? ( n284 ) : ( n341 ) ;
assign n343 =  ( n279 ) ? ( n282 ) : ( n342 ) ;
assign n344 =  ( n277 ) ? ( n280 ) : ( n343 ) ;
assign n345 =  ( n274 ) ? ( n278 ) : ( n344 ) ;
assign n346 =  { ( n338 ) , ( n345 ) }  ;
assign n347 =  { ( n331 ) , ( n346 ) }  ;
assign n348 =  { ( n324 ) , ( n347 ) }  ;
assign n349 =  { ( n317 ) , ( n348 ) }  ;
assign n350 =  { ( n310 ) , ( n349 ) }  ;
assign n351 =  { ( n303 ) , ( n350 ) }  ;
assign n352 =  { ( n296 ) , ( n351 ) }  ;
assign n353 =  { ( pre_pix ) , ( n352 ) }  ;
assign n354 =  ( n227 ) ? ( stencil_8 ) : ( n353 ) ;
assign n355 =  ( n17 ) ? ( stencil_8 ) : ( stencil_8 ) ;
assign n356 =  ( n6 ) ? ( n354 ) : ( n355 ) ;
assign n357 =  ( n4 ) ? ( stencil_8 ) : ( n356 ) ;
assign n358 = ~ ( n4 ) ;
assign n359 =  ( 1'b1 ) & ( n358 )  ;
assign n360 = ~ ( n6 ) ;
assign n361 =  ( n359 ) & ( n360 )  ;
assign n362 = ~ ( n17 ) ;
assign n363 =  ( n361 ) & ( n362 )  ;
assign n364 =  ( n361 ) & ( n17 )  ;
assign n365 =  ( n359 ) & ( n6 )  ;
assign n366 = ~ ( n23 ) ;
assign n367 =  ( n365 ) & ( n366 )  ;
assign n368 = ~ ( n274 ) ;
assign n369 =  ( n367 ) & ( n368 )  ;
assign n370 =  ( n367 ) & ( n274 )  ;
assign n371 =  ( n365 ) & ( n23 )  ;
assign n372 =  ( 1'b1 ) & ( n4 )  ;
assign RAM_0_addr0 = n370 ? (n275) : (0);
assign RAM_0_data0 = n370 ? (pre_pix) : ('dx);
assign RAM_0_wen0 = n370 ? ( 1'b1 ) : (1'b0);
assign n373 = ~ ( n277 ) ;
assign n374 =  ( n367 ) & ( n373 )  ;
assign n375 =  ( n367 ) & ( n277 )  ;
assign RAM_1_addr0 = n375 ? (n275) : (0);
assign RAM_1_data0 = n375 ? (pre_pix) : ('dx);
assign RAM_1_wen0 = n375 ? ( 1'b1 ) : (1'b0);
assign n376 = ~ ( n279 ) ;
assign n377 =  ( n367 ) & ( n376 )  ;
assign n378 =  ( n367 ) & ( n279 )  ;
assign RAM_2_addr0 = n378 ? (n275) : (0);
assign RAM_2_data0 = n378 ? (pre_pix) : ('dx);
assign RAM_2_wen0 = n378 ? ( 1'b1 ) : (1'b0);
assign n379 = ~ ( n281 ) ;
assign n380 =  ( n367 ) & ( n379 )  ;
assign n381 =  ( n367 ) & ( n281 )  ;
assign RAM_3_addr0 = n381 ? (n275) : (0);
assign RAM_3_data0 = n381 ? (pre_pix) : ('dx);
assign RAM_3_wen0 = n381 ? ( 1'b1 ) : (1'b0);
assign n382 = ~ ( n283 ) ;
assign n383 =  ( n367 ) & ( n382 )  ;
assign n384 =  ( n367 ) & ( n283 )  ;
assign RAM_4_addr0 = n384 ? (n275) : (0);
assign RAM_4_data0 = n384 ? (pre_pix) : ('dx);
assign RAM_4_wen0 = n384 ? ( 1'b1 ) : (1'b0);
assign n385 = ~ ( n285 ) ;
assign n386 =  ( n367 ) & ( n385 )  ;
assign n387 =  ( n367 ) & ( n285 )  ;
assign RAM_5_addr0 = n387 ? (n275) : (0);
assign RAM_5_data0 = n387 ? (pre_pix) : ('dx);
assign RAM_5_wen0 = n387 ? ( 1'b1 ) : (1'b0);
assign n388 = ~ ( n287 ) ;
assign n389 =  ( n367 ) & ( n388 )  ;
assign n390 =  ( n367 ) & ( n287 )  ;
assign RAM_6_addr0 = n390 ? (n275) : (0);
assign RAM_6_data0 = n390 ? (pre_pix) : ('dx);
assign RAM_6_wen0 = n390 ? ( 1'b1 ) : (1'b0);
assign n391 = ~ ( n8 ) ;
assign n392 =  ( n367 ) & ( n391 )  ;
assign n393 =  ( n367 ) & ( n8 )  ;
assign RAM_7_addr0 = n393 ? (n275) : (0);
assign RAM_7_data0 = n393 ? (pre_pix) : ('dx);
assign RAM_7_wen0 = n393 ? ( 1'b1 ) : (1'b0);
always @(posedge clk) begin
   if(rst) begin
       RAM_w <= RAM_w;
       RAM_x <= RAM_x;
       RAM_y <= RAM_y;
       arg_0_TDATA <= arg_0_TDATA;
       arg_0_TVALID <= arg_0_TVALID;
       arg_1_TREADY <= arg_1_TREADY;
       cur_pix <= cur_pix;
       gbit <= gbit;
       pre_pix <= pre_pix;
       proc_in <= proc_in;
       st_ready <= st_ready;
       stencil_0 <= stencil_0;
       stencil_1 <= stencil_1;
       stencil_2 <= stencil_2;
       stencil_3 <= stencil_3;
       stencil_4 <= stencil_4;
       stencil_5 <= stencil_5;
       stencil_6 <= stencil_6;
       stencil_7 <= stencil_7;
       stencil_8 <= stencil_8;
   end
   else if(step) begin
       RAM_w <= n20;
       RAM_x <= n29;
       RAM_y <= n36;
       arg_0_TDATA <= n214;
       arg_0_TVALID <= n220;
       arg_1_TREADY <= n232;
       cur_pix <= n235;
       gbit <= gbit;
       pre_pix <= n237;
       proc_in <= n239;
       st_ready <= n241;
       stencil_0 <= n245;
       stencil_1 <= n249;
       stencil_2 <= n253;
       stencil_3 <= n257;
       stencil_4 <= n261;
       stencil_5 <= n265;
       stencil_6 <= n269;
       stencil_7 <= n273;
       stencil_8 <= n357;
       if (RAM_0_wen0) begin
           RAM_0 [ RAM_0_addr0 ] <= RAM_0_data0 ;
       end
       if (RAM_1_wen0) begin
           RAM_1 [ RAM_1_addr0 ] <= RAM_1_data0 ;
       end
       if (RAM_2_wen0) begin
           RAM_2 [ RAM_2_addr0 ] <= RAM_2_data0 ;
       end
       if (RAM_3_wen0) begin
           RAM_3 [ RAM_3_addr0 ] <= RAM_3_data0 ;
       end
       if (RAM_4_wen0) begin
           RAM_4 [ RAM_4_addr0 ] <= RAM_4_data0 ;
       end
       if (RAM_5_wen0) begin
           RAM_5 [ RAM_5_addr0 ] <= RAM_5_data0 ;
       end
       if (RAM_6_wen0) begin
           RAM_6 [ RAM_6_addr0 ] <= RAM_6_data0 ;
       end
       if (RAM_7_wen0) begin
           RAM_7 [ RAM_7_addr0 ] <= RAM_7_data0 ;
       end
   end
end
endmodule
