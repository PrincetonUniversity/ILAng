/* PREHEADER */
module fun_gb_fun (
    input [647:0] arg1,
    output [7:0] result
);
//TODO: Add the specific function HERE.
endmodule

/* END OF PREHEADER */
module SPEC_B(
arg_0_TREADY,
arg_1_TDATA,
arg_1_TVALID,
LB1D_buff,
LB1D_in,
LB1D_it_1,
LB1D_p_cnt,
LB1D_uIn,
LB2D_proc_w,
LB2D_proc_x,
LB2D_proc_y,
LB2D_shift_0,
LB2D_shift_1,
LB2D_shift_2,
LB2D_shift_3,
LB2D_shift_4,
LB2D_shift_5,
LB2D_shift_6,
LB2D_shift_7,
LB2D_shift_x,
LB2D_shift_y,
arg_0_TDATA,
arg_0_TVALID,
arg_1_TREADY,
gb_exit_it_1,
gb_exit_it_2,
gb_exit_it_3,
gb_exit_it_4,
gb_exit_it_5,
gb_exit_it_6,
gb_exit_it_7,
gb_exit_it_8,
gb_p_cnt,
gb_pp_it_1,
gb_pp_it_2,
gb_pp_it_3,
gb_pp_it_4,
gb_pp_it_5,
gb_pp_it_6,
gb_pp_it_7,
gb_pp_it_8,
gb_pp_it_9,
in_stream_buff_0,
in_stream_buff_1,
in_stream_empty,
in_stream_full,
slice_stream_buff_0,
slice_stream_buff_1,
slice_stream_empty,
slice_stream_full,
stencil_stream_buff_0,
stencil_stream_buff_1,
stencil_stream_empty,
stencil_stream_full,
clk,rst,
step
);
input            arg_0_TREADY;
input      [7:0] arg_1_TDATA;
input            arg_1_TVALID;
input clk;
input rst;
input step;
output      [7:0] LB1D_buff;
output      [7:0] LB1D_in;
output            LB1D_it_1;
output     [18:0] LB1D_p_cnt;
output      [7:0] LB1D_uIn;
output     [63:0] LB2D_proc_w;
output      [8:0] LB2D_proc_x;
output      [9:0] LB2D_proc_y;
output     [71:0] LB2D_shift_0;
output     [71:0] LB2D_shift_1;
output     [71:0] LB2D_shift_2;
output     [71:0] LB2D_shift_3;
output     [71:0] LB2D_shift_4;
output     [71:0] LB2D_shift_5;
output     [71:0] LB2D_shift_6;
output     [71:0] LB2D_shift_7;
output      [8:0] LB2D_shift_x;
output      [9:0] LB2D_shift_y;
output      [7:0] arg_0_TDATA;
output            arg_0_TVALID;
output            arg_1_TREADY;
output            gb_exit_it_1;
output            gb_exit_it_2;
output            gb_exit_it_3;
output            gb_exit_it_4;
output            gb_exit_it_5;
output            gb_exit_it_6;
output            gb_exit_it_7;
output            gb_exit_it_8;
output     [18:0] gb_p_cnt;
output            gb_pp_it_1;
output            gb_pp_it_2;
output            gb_pp_it_3;
output            gb_pp_it_4;
output            gb_pp_it_5;
output            gb_pp_it_6;
output            gb_pp_it_7;
output            gb_pp_it_8;
output            gb_pp_it_9;
output      [7:0] in_stream_buff_0;
output      [7:0] in_stream_buff_1;
output            in_stream_empty;
output            in_stream_full;
output     [71:0] slice_stream_buff_0;
output     [71:0] slice_stream_buff_1;
output            slice_stream_empty;
output            slice_stream_full;
output    [647:0] stencil_stream_buff_0;
output    [647:0] stencil_stream_buff_1;
output            stencil_stream_empty;
output            stencil_stream_full;
reg      [7:0] LB1D_buff;
reg      [7:0] LB1D_in;
reg            LB1D_it_1;
reg     [18:0] LB1D_p_cnt;
reg      [7:0] LB1D_uIn;
reg     [63:0] LB2D_proc_w;
reg      [8:0] LB2D_proc_x;
reg      [9:0] LB2D_proc_y;
reg     [71:0] LB2D_shift_0;
reg     [71:0] LB2D_shift_1;
reg     [71:0] LB2D_shift_2;
reg     [71:0] LB2D_shift_3;
reg     [71:0] LB2D_shift_4;
reg     [71:0] LB2D_shift_5;
reg     [71:0] LB2D_shift_6;
reg     [71:0] LB2D_shift_7;
reg      [8:0] LB2D_shift_x;
reg      [9:0] LB2D_shift_y;
reg      [7:0] arg_0_TDATA;
reg            arg_0_TVALID;
reg            arg_1_TREADY;
reg            gb_exit_it_1;
reg            gb_exit_it_2;
reg            gb_exit_it_3;
reg            gb_exit_it_4;
reg            gb_exit_it_5;
reg            gb_exit_it_6;
reg            gb_exit_it_7;
reg            gb_exit_it_8;
reg     [18:0] gb_p_cnt;
reg            gb_pp_it_1;
reg            gb_pp_it_2;
reg            gb_pp_it_3;
reg            gb_pp_it_4;
reg            gb_pp_it_5;
reg            gb_pp_it_6;
reg            gb_pp_it_7;
reg            gb_pp_it_8;
reg            gb_pp_it_9;
reg      [7:0] in_stream_buff_0;
reg      [7:0] in_stream_buff_1;
reg            in_stream_empty;
reg            in_stream_full;
reg     [71:0] slice_stream_buff_0;
reg     [71:0] slice_stream_buff_1;
reg            slice_stream_empty;
reg            slice_stream_full;
reg    [647:0] stencil_stream_buff_0;
reg    [647:0] stencil_stream_buff_1;
reg            stencil_stream_empty;
reg            stencil_stream_full;
wire            arg_0_TREADY;
wire      [7:0] arg_1_TDATA;
wire            arg_1_TVALID;
wire            n0;
wire            n1;
wire            n2;
wire            n3;
wire            n4;
wire            n5;
wire            n6;
wire            n7;
wire            n8;
wire            n9;
wire            n10;
wire            n11;
wire            n12;
wire            n13;
wire            n14;
wire            n15;
wire            n16;
wire            n17;
wire            n18;
wire            n19;
wire            n20;
wire            n21;
wire            n22;
wire            n23;
wire            n24;
wire            n25;
wire            n26;
wire            n27;
wire            n28;
wire            n29;
wire            n30;
wire            n31;
wire            n32;
wire            n33;
wire      [7:0] n34;
wire      [7:0] n35;
wire      [7:0] n36;
wire      [7:0] n37;
wire      [7:0] n38;
wire      [7:0] n39;
wire      [7:0] n40;
wire      [7:0] n41;
wire      [7:0] n42;
wire      [7:0] n43;
wire      [7:0] n44;
wire      [7:0] n45;
wire            n46;
wire            n47;
wire            n48;
wire            n49;
wire            n50;
wire     [18:0] n51;
wire     [18:0] n52;
wire     [18:0] n53;
wire     [18:0] n54;
wire     [18:0] n55;
wire     [18:0] n56;
wire     [18:0] n57;
wire     [18:0] n58;
wire      [7:0] n59;
wire      [7:0] n60;
wire      [7:0] n61;
wire      [7:0] n62;
wire      [7:0] n63;
wire            n64;
wire            n65;
wire     [63:0] n66;
wire     [63:0] n67;
wire     [63:0] n68;
wire     [63:0] n69;
wire     [63:0] n70;
wire     [63:0] n71;
wire     [63:0] n72;
wire     [63:0] n73;
wire     [63:0] n74;
wire      [8:0] n75;
wire      [8:0] n76;
wire      [8:0] n77;
wire      [8:0] n78;
wire      [8:0] n79;
wire      [8:0] n80;
wire      [8:0] n81;
wire      [8:0] n82;
wire            n83;
wire      [9:0] n84;
wire      [9:0] n85;
wire      [9:0] n86;
wire      [9:0] n87;
wire      [9:0] n88;
wire      [9:0] n89;
wire      [9:0] n90;
wire      [9:0] n91;
wire      [9:0] n92;
wire     [71:0] n93;
wire     [71:0] n94;
wire     [71:0] n95;
wire     [71:0] n96;
wire     [71:0] n97;
wire     [71:0] n98;
wire     [71:0] n99;
wire     [71:0] n100;
wire     [71:0] n101;
wire     [71:0] n102;
wire     [71:0] n103;
wire     [71:0] n104;
wire     [71:0] n105;
wire     [71:0] n106;
wire     [71:0] n107;
wire     [71:0] n108;
wire     [71:0] n109;
wire     [71:0] n110;
wire     [71:0] n111;
wire     [71:0] n112;
wire     [71:0] n113;
wire     [71:0] n114;
wire     [71:0] n115;
wire     [71:0] n116;
wire     [71:0] n117;
wire     [71:0] n118;
wire     [71:0] n119;
wire     [71:0] n120;
wire     [71:0] n121;
wire     [71:0] n122;
wire     [71:0] n123;
wire     [71:0] n124;
wire     [71:0] n125;
wire     [71:0] n126;
wire     [71:0] n127;
wire     [71:0] n128;
wire     [71:0] n129;
wire     [71:0] n130;
wire     [71:0] n131;
wire     [71:0] n132;
wire     [71:0] n133;
wire     [71:0] n134;
wire            n135;
wire     [71:0] n136;
wire     [71:0] n137;
wire     [71:0] n138;
wire     [71:0] n139;
wire     [71:0] n140;
wire     [71:0] n141;
wire     [71:0] n142;
wire            n143;
wire      [8:0] n144;
wire      [8:0] n145;
wire      [8:0] n146;
wire      [8:0] n147;
wire      [8:0] n148;
wire      [8:0] n149;
wire      [8:0] n150;
wire      [8:0] n151;
wire            n152;
wire            n153;
wire      [9:0] n154;
wire      [9:0] n155;
wire      [9:0] n156;
wire      [9:0] n157;
wire      [9:0] n158;
wire      [9:0] n159;
wire      [9:0] n160;
wire      [9:0] n161;
wire      [9:0] n162;
wire            n163;
wire    [647:0] n164;
wire      [7:0] n165;
wire      [7:0] n167;
wire      [7:0] n168;
wire      [7:0] n169;
wire      [7:0] n170;
wire      [7:0] n171;
wire      [7:0] n172;
wire      [7:0] n173;
wire            n174;
wire            n175;
wire            n176;
wire            n177;
wire            n178;
wire            n179;
wire            n180;
wire            n181;
wire            n182;
wire            n183;
wire            n184;
wire            n185;
wire            n186;
wire            n187;
wire            n188;
wire            n189;
wire            n190;
wire            n191;
wire            n192;
wire            n193;
wire            n194;
wire            n195;
wire            n196;
wire            n197;
wire            n198;
wire            n199;
wire            n200;
wire            n201;
wire            n202;
wire            n203;
wire            n204;
wire            n205;
wire            n206;
wire            n207;
wire            n208;
wire            n209;
wire            n210;
wire            n211;
wire            n212;
wire            n213;
wire            n214;
wire            n215;
wire            n216;
wire            n217;
wire            n218;
wire            n219;
wire            n220;
wire            n221;
wire            n222;
wire            n223;
wire            n224;
wire            n225;
wire            n226;
wire            n227;
wire            n228;
wire            n229;
wire            n230;
wire            n231;
wire            n232;
wire            n233;
wire            n234;
wire            n235;
wire            n236;
wire            n237;
wire            n238;
wire            n239;
wire            n240;
wire     [18:0] n241;
wire     [18:0] n242;
wire     [18:0] n243;
wire     [18:0] n244;
wire     [18:0] n245;
wire     [18:0] n246;
wire     [18:0] n247;
wire     [18:0] n248;
wire            n249;
wire            n250;
wire            n251;
wire            n252;
wire            n253;
wire            n254;
wire            n255;
wire            n256;
wire            n257;
wire            n258;
wire            n259;
wire            n260;
wire            n261;
wire            n262;
wire            n263;
wire            n264;
wire            n265;
wire            n266;
wire            n267;
wire            n268;
wire            n269;
wire            n270;
wire            n271;
wire            n272;
wire            n273;
wire            n274;
wire            n275;
wire            n276;
wire            n277;
wire            n278;
wire            n279;
wire            n280;
wire            n281;
wire            n282;
wire            n283;
wire            n284;
wire            n285;
wire            n286;
wire            n287;
wire            n288;
wire            n289;
wire            n290;
wire            n291;
wire            n292;
wire            n293;
wire            n294;
wire            n295;
wire            n296;
wire            n297;
wire            n298;
wire            n299;
wire            n300;
wire            n301;
wire            n302;
wire      [7:0] n303;
wire      [7:0] n304;
wire      [7:0] n305;
wire      [7:0] n306;
wire      [7:0] n307;
wire      [7:0] n308;
wire      [7:0] n309;
wire      [7:0] n310;
wire      [7:0] n311;
wire      [7:0] n312;
wire      [7:0] n313;
wire      [7:0] n314;
wire            n315;
wire            n316;
wire            n317;
wire            n318;
wire            n319;
wire            n320;
wire            n321;
wire            n322;
wire            n323;
wire            n324;
wire            n325;
wire            n326;
wire            n327;
wire            n328;
wire            n329;
wire            n330;
wire      [7:0] n331;
wire            n332;
wire      [8:0] n333;
wire      [7:0] n334;
wire            n335;
wire      [7:0] n336;
wire            n337;
wire      [7:0] n338;
wire            n339;
wire      [7:0] n340;
wire            n341;
wire      [7:0] n342;
wire            n343;
wire      [7:0] n344;
wire            n345;
wire      [7:0] n346;
wire      [7:0] n347;
wire      [7:0] n348;
wire      [7:0] n349;
wire      [7:0] n350;
wire      [7:0] n351;
wire      [7:0] n352;
wire      [7:0] n353;
wire      [7:0] n354;
wire      [7:0] n355;
wire      [7:0] n356;
wire      [7:0] n357;
wire      [7:0] n358;
wire      [7:0] n359;
wire      [7:0] n360;
wire      [7:0] n361;
wire      [7:0] n362;
wire      [7:0] n363;
wire      [7:0] n364;
wire      [7:0] n365;
wire      [7:0] n366;
wire      [7:0] n367;
wire      [7:0] n368;
wire      [7:0] n369;
wire      [7:0] n370;
wire      [7:0] n371;
wire      [7:0] n372;
wire      [7:0] n373;
wire      [7:0] n374;
wire      [7:0] n375;
wire      [7:0] n376;
wire      [7:0] n377;
wire      [7:0] n378;
wire      [7:0] n379;
wire      [7:0] n380;
wire      [7:0] n381;
wire      [7:0] n382;
wire      [7:0] n383;
wire      [7:0] n384;
wire      [7:0] n385;
wire      [7:0] n386;
wire      [7:0] n387;
wire      [7:0] n388;
wire      [7:0] n389;
wire      [7:0] n390;
wire      [7:0] n391;
wire      [7:0] n392;
wire      [7:0] n393;
wire      [7:0] n394;
wire      [7:0] n395;
wire      [7:0] n396;
wire      [7:0] n397;
wire      [7:0] n398;
wire      [7:0] n399;
wire      [7:0] n400;
wire      [7:0] n401;
wire      [7:0] n402;
wire      [7:0] n403;
wire     [15:0] n404;
wire     [23:0] n405;
wire     [31:0] n406;
wire     [39:0] n407;
wire     [47:0] n408;
wire     [55:0] n409;
wire     [63:0] n410;
wire     [71:0] n411;
wire     [71:0] n412;
wire     [71:0] n413;
wire     [71:0] n414;
wire     [71:0] n415;
wire     [71:0] n416;
wire     [71:0] n417;
wire     [71:0] n418;
wire     [71:0] n419;
wire     [71:0] n420;
wire     [71:0] n421;
wire     [71:0] n422;
wire     [71:0] n423;
wire     [71:0] n424;
wire     [71:0] n425;
wire            n426;
wire            n427;
wire            n428;
wire            n429;
wire            n430;
wire            n431;
wire            n432;
wire            n433;
wire            n434;
wire            n435;
wire            n436;
wire            n437;
wire            n438;
wire            n439;
wire            n440;
wire            n441;
wire            n442;
wire            n443;
wire            n444;
wire            n445;
wire      [7:0] n446;
wire      [7:0] n447;
wire      [7:0] n448;
wire      [7:0] n449;
wire      [7:0] n450;
wire      [7:0] n451;
wire      [7:0] n452;
wire      [7:0] n453;
wire      [7:0] n454;
wire     [15:0] n455;
wire     [23:0] n456;
wire     [31:0] n457;
wire     [39:0] n458;
wire     [47:0] n459;
wire     [55:0] n460;
wire     [63:0] n461;
wire     [71:0] n462;
wire      [7:0] n463;
wire      [7:0] n464;
wire      [7:0] n465;
wire      [7:0] n466;
wire      [7:0] n467;
wire      [7:0] n468;
wire      [7:0] n469;
wire      [7:0] n470;
wire      [7:0] n471;
wire     [15:0] n472;
wire     [23:0] n473;
wire     [31:0] n474;
wire     [39:0] n475;
wire     [47:0] n476;
wire     [55:0] n477;
wire     [63:0] n478;
wire     [71:0] n479;
wire      [7:0] n480;
wire      [7:0] n481;
wire      [7:0] n482;
wire      [7:0] n483;
wire      [7:0] n484;
wire      [7:0] n485;
wire      [7:0] n486;
wire      [7:0] n487;
wire      [7:0] n488;
wire     [15:0] n489;
wire     [23:0] n490;
wire     [31:0] n491;
wire     [39:0] n492;
wire     [47:0] n493;
wire     [55:0] n494;
wire     [63:0] n495;
wire     [71:0] n496;
wire      [7:0] n497;
wire      [7:0] n498;
wire      [7:0] n499;
wire      [7:0] n500;
wire      [7:0] n501;
wire      [7:0] n502;
wire      [7:0] n503;
wire      [7:0] n504;
wire      [7:0] n505;
wire     [15:0] n506;
wire     [23:0] n507;
wire     [31:0] n508;
wire     [39:0] n509;
wire     [47:0] n510;
wire     [55:0] n511;
wire     [63:0] n512;
wire     [71:0] n513;
wire      [7:0] n514;
wire      [7:0] n515;
wire      [7:0] n516;
wire      [7:0] n517;
wire      [7:0] n518;
wire      [7:0] n519;
wire      [7:0] n520;
wire      [7:0] n521;
wire      [7:0] n522;
wire     [15:0] n523;
wire     [23:0] n524;
wire     [31:0] n525;
wire     [39:0] n526;
wire     [47:0] n527;
wire     [55:0] n528;
wire     [63:0] n529;
wire     [71:0] n530;
wire      [7:0] n531;
wire      [7:0] n532;
wire      [7:0] n533;
wire      [7:0] n534;
wire      [7:0] n535;
wire      [7:0] n536;
wire      [7:0] n537;
wire      [7:0] n538;
wire      [7:0] n539;
wire     [15:0] n540;
wire     [23:0] n541;
wire     [31:0] n542;
wire     [39:0] n543;
wire     [47:0] n544;
wire     [55:0] n545;
wire     [63:0] n546;
wire     [71:0] n547;
wire      [7:0] n548;
wire      [7:0] n549;
wire      [7:0] n550;
wire      [7:0] n551;
wire      [7:0] n552;
wire      [7:0] n553;
wire      [7:0] n554;
wire      [7:0] n555;
wire      [7:0] n556;
wire     [15:0] n557;
wire     [23:0] n558;
wire     [31:0] n559;
wire     [39:0] n560;
wire     [47:0] n561;
wire     [55:0] n562;
wire     [63:0] n563;
wire     [71:0] n564;
wire      [7:0] n565;
wire      [7:0] n566;
wire      [7:0] n567;
wire      [7:0] n568;
wire      [7:0] n569;
wire      [7:0] n570;
wire      [7:0] n571;
wire      [7:0] n572;
wire      [7:0] n573;
wire     [15:0] n574;
wire     [23:0] n575;
wire     [31:0] n576;
wire     [39:0] n577;
wire     [47:0] n578;
wire     [55:0] n579;
wire     [63:0] n580;
wire     [71:0] n581;
wire      [7:0] n582;
wire      [7:0] n583;
wire      [7:0] n584;
wire      [7:0] n585;
wire      [7:0] n586;
wire      [7:0] n587;
wire      [7:0] n588;
wire      [7:0] n589;
wire      [7:0] n590;
wire     [15:0] n591;
wire     [23:0] n592;
wire     [31:0] n593;
wire     [39:0] n594;
wire     [47:0] n595;
wire     [55:0] n596;
wire     [63:0] n597;
wire     [71:0] n598;
wire    [143:0] n599;
wire    [215:0] n600;
wire    [287:0] n601;
wire    [359:0] n602;
wire    [431:0] n603;
wire    [503:0] n604;
wire    [575:0] n605;
wire    [647:0] n606;
wire    [647:0] n607;
wire    [647:0] n608;
wire    [647:0] n609;
wire    [647:0] n610;
wire    [647:0] n611;
wire    [647:0] n612;
wire    [647:0] n613;
wire            n614;
wire    [647:0] n615;
wire    [647:0] n616;
wire    [647:0] n617;
wire    [647:0] n618;
wire    [647:0] n619;
wire    [647:0] n620;
wire            n621;
wire            n622;
wire            n623;
wire            n624;
wire            n625;
wire            n626;
wire            n627;
wire            n628;
wire            n629;
wire            n630;
wire            n631;
wire            n632;
wire            n633;
wire            n634;
wire            n635;
wire            n636;
wire            n637;
wire            n638;
wire            n639;
wire      [8:0] LB2D_proc_0_addr0;
wire      [7:0] LB2D_proc_0_data0;
wire            LB2D_proc_0_wen0;
wire            n640;
wire            n641;
wire            n642;
wire            n643;
wire            n644;
wire            n645;
wire            n646;
wire            n647;
wire            n648;
wire            n649;
wire            n650;
wire            n651;
wire            n652;
wire            n653;
wire            n654;
wire            n655;
wire            n656;
wire            n657;
wire            n658;
wire            n659;
wire            n660;
wire      [8:0] LB2D_proc_1_addr0;
wire      [7:0] LB2D_proc_1_data0;
wire            LB2D_proc_1_wen0;
wire            n661;
wire            n662;
wire            n663;
wire      [8:0] LB2D_proc_2_addr0;
wire      [7:0] LB2D_proc_2_data0;
wire            LB2D_proc_2_wen0;
wire            n664;
wire            n665;
wire            n666;
wire      [8:0] LB2D_proc_3_addr0;
wire      [7:0] LB2D_proc_3_data0;
wire            LB2D_proc_3_wen0;
wire            n667;
wire            n668;
wire            n669;
wire      [8:0] LB2D_proc_4_addr0;
wire      [7:0] LB2D_proc_4_data0;
wire            LB2D_proc_4_wen0;
wire            n670;
wire            n671;
wire            n672;
wire      [8:0] LB2D_proc_5_addr0;
wire      [7:0] LB2D_proc_5_data0;
wire            LB2D_proc_5_wen0;
wire            n673;
wire            n674;
wire            n675;
wire      [8:0] LB2D_proc_6_addr0;
wire      [7:0] LB2D_proc_6_data0;
wire            LB2D_proc_6_wen0;
wire            n676;
wire            n677;
wire            n678;
wire      [8:0] LB2D_proc_7_addr0;
wire      [7:0] LB2D_proc_7_data0;
wire            LB2D_proc_7_wen0;
wire            n679;
wire            n680;
wire            n681;
reg      [7:0] LB2D_proc_0[511:0];
reg      [7:0] LB2D_proc_1[511:0];
reg      [7:0] LB2D_proc_2[511:0];
reg      [7:0] LB2D_proc_3[511:0];
reg      [7:0] LB2D_proc_4[511:0];
reg      [7:0] LB2D_proc_5[511:0];
reg      [7:0] LB2D_proc_6[511:0];
reg      [7:0] LB2D_proc_7[511:0];
wire clk;
wire rst;
wire step;
assign n0 =  ( arg_0_TREADY ) == ( 1'd1 )  ;
assign n1 =  ( arg_0_TVALID ) == ( 1'd1 )  ;
assign n2 =  ( n0 ) & ( n1 )  ;
assign n3 =  ( arg_1_TVALID ) == ( 1'd0 )  ;
assign n4 =  ( n2 ) & ( n3 )  ;
assign n5 =  ( arg_1_TREADY ) == ( 1'd1 )  ;
assign n6 =  ( arg_1_TVALID ) == ( 1'd1 )  ;
assign n7 =  ( n5 ) & ( n6 )  ;
assign n8 =  ( arg_0_TREADY ) == ( 1'd0 )  ;
assign n9 =  ( n7 ) & ( n8 )  ;
assign n10 =  ( arg_0_TVALID ) == ( 1'd0 )  ;
assign n11 =  ( gb_exit_it_1 ) == ( 1'd0 )  ;
assign n12 =  ( stencil_stream_empty ) == ( 1'd0 )  ;
assign n13 =  ( n11 ) & ( n12 )  ;
assign n14 =  ( gb_exit_it_1 ) == ( 1'd1 )  ;
assign n15 =  ( gb_exit_it_8 ) == ( 1'd0 )  ;
assign n16 =  ( n14 ) & ( n15 )  ;
assign n17 =  ( n13 ) | ( n16 )  ;
assign n18 =  ( n10 ) & ( n17 )  ;
assign n19 =  ( slice_stream_empty ) == ( 1'd0 )  ;
assign n20 =  ( stencil_stream_full ) == ( 1'd0 )  ;
assign n21 =  ( LB2D_shift_x ) < ( 9'd8 )  ;
assign n22 =  ( LB2D_shift_x ) > ( 9'd0 )  ;
assign n23 =  ( n21 ) & ( n22 )  ;
assign n24 =  ( n20 ) | ( n23 )  ;
assign n25 =  ( n19 ) & ( n24 )  ;
assign n26 =  ( in_stream_empty ) == ( 1'd0 )  ;
assign n27 =  ( slice_stream_full ) == ( 1'd0 )  ;
assign n28 =  ( LB2D_proc_y ) < ( 10'd8 )  ;
assign n29 =  ( n27 ) | ( n28 )  ;
assign n30 =  ( n26 ) & ( n29 )  ;
assign n31 =  ( arg_1_TREADY ) == ( 1'd0 )  ;
assign n32 =  ( in_stream_full ) == ( 1'd0 )  ;
assign n33 =  ( n31 ) & ( n32 )  ;
assign n34 =  ( n33 ) ? ( LB1D_uIn ) : ( LB1D_buff ) ;
assign n35 =  ( n30 ) ? ( LB1D_buff ) : ( n34 ) ;
assign n36 =  ( n25 ) ? ( LB1D_buff ) : ( n35 ) ;
assign n37 =  ( n18 ) ? ( LB1D_buff ) : ( n36 ) ;
assign n38 =  ( n9 ) ? ( LB1D_buff ) : ( n37 ) ;
assign n39 =  ( n4 ) ? ( LB1D_buff ) : ( n38 ) ;
assign n40 =  ( n33 ) ? ( LB1D_in ) : ( LB1D_in ) ;
assign n41 =  ( n30 ) ? ( LB1D_in ) : ( n40 ) ;
assign n42 =  ( n25 ) ? ( LB1D_in ) : ( n41 ) ;
assign n43 =  ( n18 ) ? ( LB1D_in ) : ( n42 ) ;
assign n44 =  ( n9 ) ? ( arg_1_TDATA ) : ( n43 ) ;
assign n45 =  ( n4 ) ? ( LB1D_in ) : ( n44 ) ;
assign n46 =  ( LB1D_it_1 ) == ( 1'd1 )  ;
assign n47 =  ( LB1D_p_cnt ) == ( 19'd316224 )  ;
assign n48 =  ( n46 ) & ( n47 )  ;
assign n49 =  ( n48 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n50 =  ( n33 ) ? ( n49 ) : ( LB1D_it_1 ) ;
assign n51 =  ( LB1D_p_cnt ) + ( 19'd1 )  ;
assign n52 =  ( n48 ) ? ( 19'd0 ) : ( n51 ) ;
assign n53 =  ( n33 ) ? ( n52 ) : ( LB1D_p_cnt ) ;
assign n54 =  ( n30 ) ? ( LB1D_p_cnt ) : ( n53 ) ;
assign n55 =  ( n25 ) ? ( LB1D_p_cnt ) : ( n54 ) ;
assign n56 =  ( n18 ) ? ( LB1D_p_cnt ) : ( n55 ) ;
assign n57 =  ( n9 ) ? ( LB1D_p_cnt ) : ( n56 ) ;
assign n58 =  ( n4 ) ? ( LB1D_p_cnt ) : ( n57 ) ;
assign n59 =  ( n33 ) ? ( LB1D_in ) : ( LB1D_uIn ) ;
assign n60 =  ( n30 ) ? ( LB1D_uIn ) : ( n59 ) ;
assign n61 =  ( n25 ) ? ( LB1D_uIn ) : ( n60 ) ;
assign n62 =  ( n18 ) ? ( LB1D_uIn ) : ( n61 ) ;
assign n63 =  ( n9 ) ? ( LB1D_uIn ) : ( n62 ) ;
assign n64 =  ( LB2D_proc_x ) == ( 9'd488 )  ;
assign n65 =  ( LB2D_proc_w ) == ( 64'd7 )  ;
assign n66 =  ( LB2D_proc_w ) + ( 64'd1 )  ;
assign n67 =  ( n65 ) ? ( 64'd0 ) : ( n66 ) ;
assign n68 =  ( n64 ) ? ( n67 ) : ( LB2D_proc_w ) ;
assign n69 =  ( n33 ) ? ( LB2D_proc_w ) : ( LB2D_proc_w ) ;
assign n70 =  ( n30 ) ? ( n68 ) : ( n69 ) ;
assign n71 =  ( n25 ) ? ( LB2D_proc_w ) : ( n70 ) ;
assign n72 =  ( n18 ) ? ( LB2D_proc_w ) : ( n71 ) ;
assign n73 =  ( n9 ) ? ( LB2D_proc_w ) : ( n72 ) ;
assign n74 =  ( n4 ) ? ( LB2D_proc_w ) : ( n73 ) ;
assign n75 =  ( LB2D_proc_x ) + ( 9'd1 )  ;
assign n76 =  ( n64 ) ? ( 9'd1 ) : ( n75 ) ;
assign n77 =  ( n33 ) ? ( LB2D_proc_x ) : ( LB2D_proc_x ) ;
assign n78 =  ( n30 ) ? ( n76 ) : ( n77 ) ;
assign n79 =  ( n25 ) ? ( LB2D_proc_x ) : ( n78 ) ;
assign n80 =  ( n18 ) ? ( LB2D_proc_x ) : ( n79 ) ;
assign n81 =  ( n9 ) ? ( LB2D_proc_x ) : ( n80 ) ;
assign n82 =  ( n4 ) ? ( LB2D_proc_x ) : ( n81 ) ;
assign n83 =  ( LB2D_proc_y ) == ( 10'd648 )  ;
assign n84 =  ( LB2D_proc_y ) + ( 10'd1 )  ;
assign n85 =  ( n83 ) ? ( 10'd0 ) : ( n84 ) ;
assign n86 =  ( n64 ) ? ( n85 ) : ( LB2D_proc_y ) ;
assign n87 =  ( n33 ) ? ( LB2D_proc_y ) : ( LB2D_proc_y ) ;
assign n88 =  ( n30 ) ? ( n86 ) : ( n87 ) ;
assign n89 =  ( n25 ) ? ( LB2D_proc_y ) : ( n88 ) ;
assign n90 =  ( n18 ) ? ( LB2D_proc_y ) : ( n89 ) ;
assign n91 =  ( n9 ) ? ( LB2D_proc_y ) : ( n90 ) ;
assign n92 =  ( n4 ) ? ( LB2D_proc_y ) : ( n91 ) ;
assign n93 =  ( n33 ) ? ( LB2D_shift_0 ) : ( LB2D_shift_0 ) ;
assign n94 =  ( n30 ) ? ( LB2D_shift_0 ) : ( n93 ) ;
assign n95 =  ( n25 ) ? ( LB2D_shift_1 ) : ( n94 ) ;
assign n96 =  ( n18 ) ? ( LB2D_shift_0 ) : ( n95 ) ;
assign n97 =  ( n9 ) ? ( LB2D_shift_0 ) : ( n96 ) ;
assign n98 =  ( n4 ) ? ( LB2D_shift_0 ) : ( n97 ) ;
assign n99 =  ( n33 ) ? ( LB2D_shift_1 ) : ( LB2D_shift_1 ) ;
assign n100 =  ( n30 ) ? ( LB2D_shift_1 ) : ( n99 ) ;
assign n101 =  ( n25 ) ? ( LB2D_shift_2 ) : ( n100 ) ;
assign n102 =  ( n18 ) ? ( LB2D_shift_1 ) : ( n101 ) ;
assign n103 =  ( n9 ) ? ( LB2D_shift_1 ) : ( n102 ) ;
assign n104 =  ( n4 ) ? ( LB2D_shift_1 ) : ( n103 ) ;
assign n105 =  ( n33 ) ? ( LB2D_shift_2 ) : ( LB2D_shift_2 ) ;
assign n106 =  ( n30 ) ? ( LB2D_shift_2 ) : ( n105 ) ;
assign n107 =  ( n25 ) ? ( LB2D_shift_3 ) : ( n106 ) ;
assign n108 =  ( n18 ) ? ( LB2D_shift_2 ) : ( n107 ) ;
assign n109 =  ( n9 ) ? ( LB2D_shift_2 ) : ( n108 ) ;
assign n110 =  ( n4 ) ? ( LB2D_shift_2 ) : ( n109 ) ;
assign n111 =  ( n33 ) ? ( LB2D_shift_3 ) : ( LB2D_shift_3 ) ;
assign n112 =  ( n30 ) ? ( LB2D_shift_3 ) : ( n111 ) ;
assign n113 =  ( n25 ) ? ( LB2D_shift_4 ) : ( n112 ) ;
assign n114 =  ( n18 ) ? ( LB2D_shift_3 ) : ( n113 ) ;
assign n115 =  ( n9 ) ? ( LB2D_shift_3 ) : ( n114 ) ;
assign n116 =  ( n4 ) ? ( LB2D_shift_3 ) : ( n115 ) ;
assign n117 =  ( n33 ) ? ( LB2D_shift_4 ) : ( LB2D_shift_4 ) ;
assign n118 =  ( n30 ) ? ( LB2D_shift_4 ) : ( n117 ) ;
assign n119 =  ( n25 ) ? ( LB2D_shift_5 ) : ( n118 ) ;
assign n120 =  ( n18 ) ? ( LB2D_shift_4 ) : ( n119 ) ;
assign n121 =  ( n9 ) ? ( LB2D_shift_4 ) : ( n120 ) ;
assign n122 =  ( n4 ) ? ( LB2D_shift_4 ) : ( n121 ) ;
assign n123 =  ( n33 ) ? ( LB2D_shift_5 ) : ( LB2D_shift_5 ) ;
assign n124 =  ( n30 ) ? ( LB2D_shift_5 ) : ( n123 ) ;
assign n125 =  ( n25 ) ? ( LB2D_shift_6 ) : ( n124 ) ;
assign n126 =  ( n18 ) ? ( LB2D_shift_5 ) : ( n125 ) ;
assign n127 =  ( n9 ) ? ( LB2D_shift_5 ) : ( n126 ) ;
assign n128 =  ( n4 ) ? ( LB2D_shift_5 ) : ( n127 ) ;
assign n129 =  ( n33 ) ? ( LB2D_shift_6 ) : ( LB2D_shift_6 ) ;
assign n130 =  ( n30 ) ? ( LB2D_shift_6 ) : ( n129 ) ;
assign n131 =  ( n25 ) ? ( LB2D_shift_7 ) : ( n130 ) ;
assign n132 =  ( n18 ) ? ( LB2D_shift_6 ) : ( n131 ) ;
assign n133 =  ( n9 ) ? ( LB2D_shift_6 ) : ( n132 ) ;
assign n134 =  ( n4 ) ? ( LB2D_shift_6 ) : ( n133 ) ;
assign n135 =  ( slice_stream_full ) == ( 1'd1 )  ;
assign n136 =  ( n135 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n137 =  ( n33 ) ? ( LB2D_shift_7 ) : ( LB2D_shift_7 ) ;
assign n138 =  ( n30 ) ? ( LB2D_shift_7 ) : ( n137 ) ;
assign n139 =  ( n25 ) ? ( n136 ) : ( n138 ) ;
assign n140 =  ( n18 ) ? ( LB2D_shift_7 ) : ( n139 ) ;
assign n141 =  ( n9 ) ? ( LB2D_shift_7 ) : ( n140 ) ;
assign n142 =  ( n4 ) ? ( LB2D_shift_7 ) : ( n141 ) ;
assign n143 =  ( LB2D_shift_x ) == ( 9'd488 )  ;
assign n144 =  ( LB2D_shift_x ) + ( 9'd1 )  ;
assign n145 =  ( n143 ) ? ( 9'd0 ) : ( n144 ) ;
assign n146 =  ( n33 ) ? ( LB2D_shift_x ) : ( LB2D_shift_x ) ;
assign n147 =  ( n30 ) ? ( LB2D_shift_x ) : ( n146 ) ;
assign n148 =  ( n25 ) ? ( n145 ) : ( n147 ) ;
assign n149 =  ( n18 ) ? ( LB2D_shift_x ) : ( n148 ) ;
assign n150 =  ( n9 ) ? ( LB2D_shift_x ) : ( n149 ) ;
assign n151 =  ( n4 ) ? ( LB2D_shift_x ) : ( n150 ) ;
assign n152 =  ( LB2D_shift_y ) < ( 10'd640 )  ;
assign n153 =  ( LB2D_shift_x ) < ( 9'd488 )  ;
assign n154 =  ( LB2D_shift_y ) + ( 10'd1 )  ;
assign n155 =  ( n153 ) ? ( LB2D_shift_y ) : ( n154 ) ;
assign n156 =  ( n152 ) ? ( n155 ) : ( 10'd640 ) ;
assign n157 =  ( n33 ) ? ( LB2D_shift_y ) : ( LB2D_shift_y ) ;
assign n158 =  ( n30 ) ? ( LB2D_shift_y ) : ( n157 ) ;
assign n159 =  ( n25 ) ? ( n156 ) : ( n158 ) ;
assign n160 =  ( n18 ) ? ( LB2D_shift_y ) : ( n159 ) ;
assign n161 =  ( n9 ) ? ( LB2D_shift_y ) : ( n160 ) ;
assign n162 =  ( n4 ) ? ( LB2D_shift_y ) : ( n161 ) ;
assign n163 =  ( stencil_stream_full ) == ( 1'd1 )  ;
assign n164 =  ( n163 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_0 ) ;
fun_gb_fun  applyFunc_n166(
    .arg1( n164 ),
    .result( n165 )
);
assign n167 = n165 ;
assign n168 =  ( n33 ) ? ( arg_0_TDATA ) : ( arg_0_TDATA ) ;
assign n169 =  ( n30 ) ? ( arg_0_TDATA ) : ( n168 ) ;
assign n170 =  ( n25 ) ? ( arg_0_TDATA ) : ( n169 ) ;
assign n171 =  ( n18 ) ? ( n167 ) : ( n170 ) ;
assign n172 =  ( n9 ) ? ( arg_0_TDATA ) : ( n171 ) ;
assign n173 =  ( n4 ) ? ( arg_0_TDATA ) : ( n172 ) ;
assign n174 =  ( gb_pp_it_8 ) == ( 1'd1 )  ;
assign n175 =  ( gb_exit_it_7 ) == ( 1'd0 )  ;
assign n176 =  ( n174 ) & ( n175 )  ;
assign n177 =  ( n176 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n178 =  ( n33 ) ? ( arg_0_TVALID ) : ( arg_0_TVALID ) ;
assign n179 =  ( n30 ) ? ( arg_0_TVALID ) : ( n178 ) ;
assign n180 =  ( n25 ) ? ( arg_0_TVALID ) : ( n179 ) ;
assign n181 =  ( n18 ) ? ( n177 ) : ( n180 ) ;
assign n182 =  ( n9 ) ? ( arg_0_TVALID ) : ( n181 ) ;
assign n183 =  ( n4 ) ? ( 1'd0 ) : ( n182 ) ;
assign n184 =  ( n33 ) ? ( 1'd1 ) : ( arg_1_TREADY ) ;
assign n185 =  ( n30 ) ? ( arg_1_TREADY ) : ( n184 ) ;
assign n186 =  ( n25 ) ? ( arg_1_TREADY ) : ( n185 ) ;
assign n187 =  ( n18 ) ? ( arg_1_TREADY ) : ( n186 ) ;
assign n188 =  ( n9 ) ? ( 1'd0 ) : ( n187 ) ;
assign n189 =  ( n4 ) ? ( arg_1_TREADY ) : ( n188 ) ;
assign n190 =  ( gb_p_cnt ) == ( 19'd307200 )  ;
assign n191 =  ( n190 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n192 =  ( n33 ) ? ( gb_exit_it_1 ) : ( gb_exit_it_1 ) ;
assign n193 =  ( n30 ) ? ( gb_exit_it_1 ) : ( n192 ) ;
assign n194 =  ( n25 ) ? ( gb_exit_it_1 ) : ( n193 ) ;
assign n195 =  ( n18 ) ? ( n191 ) : ( n194 ) ;
assign n196 =  ( n9 ) ? ( gb_exit_it_1 ) : ( n195 ) ;
assign n197 =  ( n4 ) ? ( gb_exit_it_1 ) : ( n196 ) ;
assign n198 =  ( n33 ) ? ( gb_exit_it_2 ) : ( gb_exit_it_2 ) ;
assign n199 =  ( n30 ) ? ( gb_exit_it_2 ) : ( n198 ) ;
assign n200 =  ( n25 ) ? ( gb_exit_it_2 ) : ( n199 ) ;
assign n201 =  ( n18 ) ? ( gb_exit_it_1 ) : ( n200 ) ;
assign n202 =  ( n9 ) ? ( gb_exit_it_2 ) : ( n201 ) ;
assign n203 =  ( n4 ) ? ( gb_exit_it_2 ) : ( n202 ) ;
assign n204 =  ( n33 ) ? ( gb_exit_it_3 ) : ( gb_exit_it_3 ) ;
assign n205 =  ( n30 ) ? ( gb_exit_it_3 ) : ( n204 ) ;
assign n206 =  ( n25 ) ? ( gb_exit_it_3 ) : ( n205 ) ;
assign n207 =  ( n18 ) ? ( gb_exit_it_2 ) : ( n206 ) ;
assign n208 =  ( n9 ) ? ( gb_exit_it_3 ) : ( n207 ) ;
assign n209 =  ( n4 ) ? ( gb_exit_it_3 ) : ( n208 ) ;
assign n210 =  ( n33 ) ? ( gb_exit_it_4 ) : ( gb_exit_it_4 ) ;
assign n211 =  ( n30 ) ? ( gb_exit_it_4 ) : ( n210 ) ;
assign n212 =  ( n25 ) ? ( gb_exit_it_4 ) : ( n211 ) ;
assign n213 =  ( n18 ) ? ( gb_exit_it_3 ) : ( n212 ) ;
assign n214 =  ( n9 ) ? ( gb_exit_it_4 ) : ( n213 ) ;
assign n215 =  ( n4 ) ? ( gb_exit_it_4 ) : ( n214 ) ;
assign n216 =  ( n33 ) ? ( gb_exit_it_5 ) : ( gb_exit_it_5 ) ;
assign n217 =  ( n30 ) ? ( gb_exit_it_5 ) : ( n216 ) ;
assign n218 =  ( n25 ) ? ( gb_exit_it_5 ) : ( n217 ) ;
assign n219 =  ( n18 ) ? ( gb_exit_it_4 ) : ( n218 ) ;
assign n220 =  ( n9 ) ? ( gb_exit_it_5 ) : ( n219 ) ;
assign n221 =  ( n4 ) ? ( gb_exit_it_5 ) : ( n220 ) ;
assign n222 =  ( n33 ) ? ( gb_exit_it_6 ) : ( gb_exit_it_6 ) ;
assign n223 =  ( n30 ) ? ( gb_exit_it_6 ) : ( n222 ) ;
assign n224 =  ( n25 ) ? ( gb_exit_it_6 ) : ( n223 ) ;
assign n225 =  ( n18 ) ? ( gb_exit_it_5 ) : ( n224 ) ;
assign n226 =  ( n9 ) ? ( gb_exit_it_6 ) : ( n225 ) ;
assign n227 =  ( n4 ) ? ( gb_exit_it_6 ) : ( n226 ) ;
assign n228 =  ( n33 ) ? ( gb_exit_it_7 ) : ( gb_exit_it_7 ) ;
assign n229 =  ( n30 ) ? ( gb_exit_it_7 ) : ( n228 ) ;
assign n230 =  ( n25 ) ? ( gb_exit_it_7 ) : ( n229 ) ;
assign n231 =  ( n18 ) ? ( gb_exit_it_6 ) : ( n230 ) ;
assign n232 =  ( n9 ) ? ( gb_exit_it_7 ) : ( n231 ) ;
assign n233 =  ( n4 ) ? ( gb_exit_it_7 ) : ( n232 ) ;
assign n234 =  ( n33 ) ? ( gb_exit_it_8 ) : ( gb_exit_it_8 ) ;
assign n235 =  ( n30 ) ? ( gb_exit_it_8 ) : ( n234 ) ;
assign n236 =  ( n25 ) ? ( gb_exit_it_8 ) : ( n235 ) ;
assign n237 =  ( n18 ) ? ( gb_exit_it_7 ) : ( n236 ) ;
assign n238 =  ( n9 ) ? ( gb_exit_it_8 ) : ( n237 ) ;
assign n239 =  ( n4 ) ? ( gb_exit_it_8 ) : ( n238 ) ;
assign n240 =  ( gb_p_cnt ) < ( 19'd307200 )  ;
assign n241 =  ( gb_p_cnt ) + ( 19'd1 )  ;
assign n242 =  ( n240 ) ? ( n241 ) : ( 19'd307200 ) ;
assign n243 =  ( n33 ) ? ( gb_p_cnt ) : ( gb_p_cnt ) ;
assign n244 =  ( n30 ) ? ( gb_p_cnt ) : ( n243 ) ;
assign n245 =  ( n25 ) ? ( gb_p_cnt ) : ( n244 ) ;
assign n246 =  ( n18 ) ? ( n242 ) : ( n245 ) ;
assign n247 =  ( n9 ) ? ( gb_p_cnt ) : ( n246 ) ;
assign n248 =  ( n4 ) ? ( gb_p_cnt ) : ( n247 ) ;
assign n249 =  ( n33 ) ? ( gb_pp_it_1 ) : ( gb_pp_it_1 ) ;
assign n250 =  ( n30 ) ? ( gb_pp_it_1 ) : ( n249 ) ;
assign n251 =  ( n25 ) ? ( gb_pp_it_1 ) : ( n250 ) ;
assign n252 =  ( n18 ) ? ( 1'd1 ) : ( n251 ) ;
assign n253 =  ( n9 ) ? ( gb_pp_it_1 ) : ( n252 ) ;
assign n254 =  ( n4 ) ? ( gb_pp_it_1 ) : ( n253 ) ;
assign n255 =  ( n33 ) ? ( gb_pp_it_2 ) : ( gb_pp_it_2 ) ;
assign n256 =  ( n30 ) ? ( gb_pp_it_2 ) : ( n255 ) ;
assign n257 =  ( n25 ) ? ( gb_pp_it_2 ) : ( n256 ) ;
assign n258 =  ( n18 ) ? ( gb_pp_it_1 ) : ( n257 ) ;
assign n259 =  ( n9 ) ? ( gb_pp_it_2 ) : ( n258 ) ;
assign n260 =  ( n4 ) ? ( gb_pp_it_2 ) : ( n259 ) ;
assign n261 =  ( n33 ) ? ( gb_pp_it_3 ) : ( gb_pp_it_3 ) ;
assign n262 =  ( n30 ) ? ( gb_pp_it_3 ) : ( n261 ) ;
assign n263 =  ( n25 ) ? ( gb_pp_it_3 ) : ( n262 ) ;
assign n264 =  ( n18 ) ? ( gb_pp_it_2 ) : ( n263 ) ;
assign n265 =  ( n9 ) ? ( gb_pp_it_3 ) : ( n264 ) ;
assign n266 =  ( n4 ) ? ( gb_pp_it_3 ) : ( n265 ) ;
assign n267 =  ( n33 ) ? ( gb_pp_it_4 ) : ( gb_pp_it_4 ) ;
assign n268 =  ( n30 ) ? ( gb_pp_it_4 ) : ( n267 ) ;
assign n269 =  ( n25 ) ? ( gb_pp_it_4 ) : ( n268 ) ;
assign n270 =  ( n18 ) ? ( gb_pp_it_3 ) : ( n269 ) ;
assign n271 =  ( n9 ) ? ( gb_pp_it_4 ) : ( n270 ) ;
assign n272 =  ( n4 ) ? ( gb_pp_it_4 ) : ( n271 ) ;
assign n273 =  ( n33 ) ? ( gb_pp_it_5 ) : ( gb_pp_it_5 ) ;
assign n274 =  ( n30 ) ? ( gb_pp_it_5 ) : ( n273 ) ;
assign n275 =  ( n25 ) ? ( gb_pp_it_5 ) : ( n274 ) ;
assign n276 =  ( n18 ) ? ( gb_pp_it_4 ) : ( n275 ) ;
assign n277 =  ( n9 ) ? ( gb_pp_it_5 ) : ( n276 ) ;
assign n278 =  ( n4 ) ? ( gb_pp_it_5 ) : ( n277 ) ;
assign n279 =  ( n33 ) ? ( gb_pp_it_6 ) : ( gb_pp_it_6 ) ;
assign n280 =  ( n30 ) ? ( gb_pp_it_6 ) : ( n279 ) ;
assign n281 =  ( n25 ) ? ( gb_pp_it_6 ) : ( n280 ) ;
assign n282 =  ( n18 ) ? ( gb_pp_it_5 ) : ( n281 ) ;
assign n283 =  ( n9 ) ? ( gb_pp_it_6 ) : ( n282 ) ;
assign n284 =  ( n4 ) ? ( gb_pp_it_6 ) : ( n283 ) ;
assign n285 =  ( n33 ) ? ( gb_pp_it_7 ) : ( gb_pp_it_7 ) ;
assign n286 =  ( n30 ) ? ( gb_pp_it_7 ) : ( n285 ) ;
assign n287 =  ( n25 ) ? ( gb_pp_it_7 ) : ( n286 ) ;
assign n288 =  ( n18 ) ? ( gb_pp_it_6 ) : ( n287 ) ;
assign n289 =  ( n9 ) ? ( gb_pp_it_7 ) : ( n288 ) ;
assign n290 =  ( n4 ) ? ( gb_pp_it_7 ) : ( n289 ) ;
assign n291 =  ( n33 ) ? ( gb_pp_it_8 ) : ( gb_pp_it_8 ) ;
assign n292 =  ( n30 ) ? ( gb_pp_it_8 ) : ( n291 ) ;
assign n293 =  ( n25 ) ? ( gb_pp_it_8 ) : ( n292 ) ;
assign n294 =  ( n18 ) ? ( gb_pp_it_7 ) : ( n293 ) ;
assign n295 =  ( n9 ) ? ( gb_pp_it_8 ) : ( n294 ) ;
assign n296 =  ( n4 ) ? ( gb_pp_it_8 ) : ( n295 ) ;
assign n297 =  ( n33 ) ? ( gb_pp_it_9 ) : ( gb_pp_it_9 ) ;
assign n298 =  ( n30 ) ? ( gb_pp_it_9 ) : ( n297 ) ;
assign n299 =  ( n25 ) ? ( gb_pp_it_9 ) : ( n298 ) ;
assign n300 =  ( n18 ) ? ( gb_pp_it_8 ) : ( n299 ) ;
assign n301 =  ( n9 ) ? ( gb_pp_it_9 ) : ( n300 ) ;
assign n302 =  ( n4 ) ? ( gb_pp_it_9 ) : ( n301 ) ;
assign n303 =  ( n33 ) ? ( LB1D_uIn ) : ( in_stream_buff_0 ) ;
assign n304 =  ( n30 ) ? ( in_stream_buff_0 ) : ( n303 ) ;
assign n305 =  ( n25 ) ? ( in_stream_buff_0 ) : ( n304 ) ;
assign n306 =  ( n18 ) ? ( in_stream_buff_0 ) : ( n305 ) ;
assign n307 =  ( n9 ) ? ( in_stream_buff_0 ) : ( n306 ) ;
assign n308 =  ( n4 ) ? ( in_stream_buff_0 ) : ( n307 ) ;
assign n309 =  ( n33 ) ? ( in_stream_buff_0 ) : ( in_stream_buff_1 ) ;
assign n310 =  ( n30 ) ? ( in_stream_buff_1 ) : ( n309 ) ;
assign n311 =  ( n25 ) ? ( in_stream_buff_1 ) : ( n310 ) ;
assign n312 =  ( n18 ) ? ( in_stream_buff_1 ) : ( n311 ) ;
assign n313 =  ( n9 ) ? ( in_stream_buff_1 ) : ( n312 ) ;
assign n314 =  ( n4 ) ? ( in_stream_buff_1 ) : ( n313 ) ;
assign n315 =  ( in_stream_full ) == ( 1'd1 )  ;
assign n316 =  ( n315 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n317 =  ( n33 ) ? ( 1'd0 ) : ( in_stream_empty ) ;
assign n318 =  ( n30 ) ? ( n316 ) : ( n317 ) ;
assign n319 =  ( n25 ) ? ( in_stream_empty ) : ( n318 ) ;
assign n320 =  ( n18 ) ? ( in_stream_empty ) : ( n319 ) ;
assign n321 =  ( n9 ) ? ( in_stream_empty ) : ( n320 ) ;
assign n322 =  ( n4 ) ? ( in_stream_empty ) : ( n321 ) ;
assign n323 =  ( in_stream_empty ) == ( 1'd1 )  ;
assign n324 =  ( n323 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n325 =  ( n33 ) ? ( n324 ) : ( in_stream_full ) ;
assign n326 =  ( n30 ) ? ( 1'd0 ) : ( n325 ) ;
assign n327 =  ( n25 ) ? ( in_stream_full ) : ( n326 ) ;
assign n328 =  ( n18 ) ? ( in_stream_full ) : ( n327 ) ;
assign n329 =  ( n9 ) ? ( in_stream_full ) : ( n328 ) ;
assign n330 =  ( n4 ) ? ( in_stream_full ) : ( n329 ) ;
assign n331 =  ( n315 ) ? ( in_stream_buff_1 ) : ( in_stream_buff_0 ) ;
assign n332 =  ( LB2D_proc_w ) == ( 64'd0 )  ;
assign n333 =  ( LB2D_proc_x ) - ( 9'd1 )  ;
assign n334 =  (  LB2D_proc_7 [ n333 ] )  ;
assign n335 =  ( LB2D_proc_w ) == ( 64'd1 )  ;
assign n336 =  (  LB2D_proc_0 [ n333 ] )  ;
assign n337 =  ( LB2D_proc_w ) == ( 64'd2 )  ;
assign n338 =  (  LB2D_proc_1 [ n333 ] )  ;
assign n339 =  ( LB2D_proc_w ) == ( 64'd3 )  ;
assign n340 =  (  LB2D_proc_2 [ n333 ] )  ;
assign n341 =  ( LB2D_proc_w ) == ( 64'd4 )  ;
assign n342 =  (  LB2D_proc_3 [ n333 ] )  ;
assign n343 =  ( LB2D_proc_w ) == ( 64'd5 )  ;
assign n344 =  (  LB2D_proc_4 [ n333 ] )  ;
assign n345 =  ( LB2D_proc_w ) == ( 64'd6 )  ;
assign n346 =  (  LB2D_proc_5 [ n333 ] )  ;
assign n347 =  (  LB2D_proc_6 [ n333 ] )  ;
assign n348 =  ( n345 ) ? ( n346 ) : ( n347 ) ;
assign n349 =  ( n343 ) ? ( n344 ) : ( n348 ) ;
assign n350 =  ( n341 ) ? ( n342 ) : ( n349 ) ;
assign n351 =  ( n339 ) ? ( n340 ) : ( n350 ) ;
assign n352 =  ( n337 ) ? ( n338 ) : ( n351 ) ;
assign n353 =  ( n335 ) ? ( n336 ) : ( n352 ) ;
assign n354 =  ( n332 ) ? ( n334 ) : ( n353 ) ;
assign n355 =  ( n345 ) ? ( n344 ) : ( n346 ) ;
assign n356 =  ( n343 ) ? ( n342 ) : ( n355 ) ;
assign n357 =  ( n341 ) ? ( n340 ) : ( n356 ) ;
assign n358 =  ( n339 ) ? ( n338 ) : ( n357 ) ;
assign n359 =  ( n337 ) ? ( n336 ) : ( n358 ) ;
assign n360 =  ( n335 ) ? ( n334 ) : ( n359 ) ;
assign n361 =  ( n332 ) ? ( n347 ) : ( n360 ) ;
assign n362 =  ( n345 ) ? ( n342 ) : ( n344 ) ;
assign n363 =  ( n343 ) ? ( n340 ) : ( n362 ) ;
assign n364 =  ( n341 ) ? ( n338 ) : ( n363 ) ;
assign n365 =  ( n339 ) ? ( n336 ) : ( n364 ) ;
assign n366 =  ( n337 ) ? ( n334 ) : ( n365 ) ;
assign n367 =  ( n335 ) ? ( n347 ) : ( n366 ) ;
assign n368 =  ( n332 ) ? ( n346 ) : ( n367 ) ;
assign n369 =  ( n345 ) ? ( n340 ) : ( n342 ) ;
assign n370 =  ( n343 ) ? ( n338 ) : ( n369 ) ;
assign n371 =  ( n341 ) ? ( n336 ) : ( n370 ) ;
assign n372 =  ( n339 ) ? ( n334 ) : ( n371 ) ;
assign n373 =  ( n337 ) ? ( n347 ) : ( n372 ) ;
assign n374 =  ( n335 ) ? ( n346 ) : ( n373 ) ;
assign n375 =  ( n332 ) ? ( n344 ) : ( n374 ) ;
assign n376 =  ( n345 ) ? ( n338 ) : ( n340 ) ;
assign n377 =  ( n343 ) ? ( n336 ) : ( n376 ) ;
assign n378 =  ( n341 ) ? ( n334 ) : ( n377 ) ;
assign n379 =  ( n339 ) ? ( n347 ) : ( n378 ) ;
assign n380 =  ( n337 ) ? ( n346 ) : ( n379 ) ;
assign n381 =  ( n335 ) ? ( n344 ) : ( n380 ) ;
assign n382 =  ( n332 ) ? ( n342 ) : ( n381 ) ;
assign n383 =  ( n345 ) ? ( n336 ) : ( n338 ) ;
assign n384 =  ( n343 ) ? ( n334 ) : ( n383 ) ;
assign n385 =  ( n341 ) ? ( n347 ) : ( n384 ) ;
assign n386 =  ( n339 ) ? ( n346 ) : ( n385 ) ;
assign n387 =  ( n337 ) ? ( n344 ) : ( n386 ) ;
assign n388 =  ( n335 ) ? ( n342 ) : ( n387 ) ;
assign n389 =  ( n332 ) ? ( n340 ) : ( n388 ) ;
assign n390 =  ( n345 ) ? ( n334 ) : ( n336 ) ;
assign n391 =  ( n343 ) ? ( n347 ) : ( n390 ) ;
assign n392 =  ( n341 ) ? ( n346 ) : ( n391 ) ;
assign n393 =  ( n339 ) ? ( n344 ) : ( n392 ) ;
assign n394 =  ( n337 ) ? ( n342 ) : ( n393 ) ;
assign n395 =  ( n335 ) ? ( n340 ) : ( n394 ) ;
assign n396 =  ( n332 ) ? ( n338 ) : ( n395 ) ;
assign n397 =  ( n345 ) ? ( n347 ) : ( n334 ) ;
assign n398 =  ( n343 ) ? ( n346 ) : ( n397 ) ;
assign n399 =  ( n341 ) ? ( n344 ) : ( n398 ) ;
assign n400 =  ( n339 ) ? ( n342 ) : ( n399 ) ;
assign n401 =  ( n337 ) ? ( n340 ) : ( n400 ) ;
assign n402 =  ( n335 ) ? ( n338 ) : ( n401 ) ;
assign n403 =  ( n332 ) ? ( n336 ) : ( n402 ) ;
assign n404 =  { ( n396 ) , ( n403 ) }  ;
assign n405 =  { ( n389 ) , ( n404 ) }  ;
assign n406 =  { ( n382 ) , ( n405 ) }  ;
assign n407 =  { ( n375 ) , ( n406 ) }  ;
assign n408 =  { ( n368 ) , ( n407 ) }  ;
assign n409 =  { ( n361 ) , ( n408 ) }  ;
assign n410 =  { ( n354 ) , ( n409 ) }  ;
assign n411 =  { ( n331 ) , ( n410 ) }  ;
assign n412 =  ( n28 ) ? ( slice_stream_buff_0 ) : ( n411 ) ;
assign n413 =  ( n33 ) ? ( slice_stream_buff_0 ) : ( slice_stream_buff_0 ) ;
assign n414 =  ( n30 ) ? ( n412 ) : ( n413 ) ;
assign n415 =  ( n25 ) ? ( slice_stream_buff_0 ) : ( n414 ) ;
assign n416 =  ( n18 ) ? ( slice_stream_buff_0 ) : ( n415 ) ;
assign n417 =  ( n9 ) ? ( slice_stream_buff_0 ) : ( n416 ) ;
assign n418 =  ( n4 ) ? ( slice_stream_buff_0 ) : ( n417 ) ;
assign n419 =  ( n28 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n420 =  ( n33 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_1 ) ;
assign n421 =  ( n30 ) ? ( n419 ) : ( n420 ) ;
assign n422 =  ( n25 ) ? ( slice_stream_buff_1 ) : ( n421 ) ;
assign n423 =  ( n18 ) ? ( slice_stream_buff_1 ) : ( n422 ) ;
assign n424 =  ( n9 ) ? ( slice_stream_buff_1 ) : ( n423 ) ;
assign n425 =  ( n4 ) ? ( slice_stream_buff_1 ) : ( n424 ) ;
assign n426 =  ( n135 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n427 =  ( n28 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n428 =  ( n33 ) ? ( slice_stream_empty ) : ( slice_stream_empty ) ;
assign n429 =  ( n30 ) ? ( n427 ) : ( n428 ) ;
assign n430 =  ( n25 ) ? ( n426 ) : ( n429 ) ;
assign n431 =  ( n18 ) ? ( slice_stream_empty ) : ( n430 ) ;
assign n432 =  ( n9 ) ? ( slice_stream_empty ) : ( n431 ) ;
assign n433 =  ( n4 ) ? ( slice_stream_empty ) : ( n432 ) ;
assign n434 =  ( slice_stream_empty ) == ( 1'd1 )  ;
assign n435 =  ( n434 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n436 =  ( n28 ) ? ( 1'd0 ) : ( n435 ) ;
assign n437 =  ( n33 ) ? ( slice_stream_full ) : ( slice_stream_full ) ;
assign n438 =  ( n30 ) ? ( n436 ) : ( n437 ) ;
assign n439 =  ( n25 ) ? ( 1'd0 ) : ( n438 ) ;
assign n440 =  ( n18 ) ? ( slice_stream_full ) : ( n439 ) ;
assign n441 =  ( n9 ) ? ( slice_stream_full ) : ( n440 ) ;
assign n442 =  ( n4 ) ? ( slice_stream_full ) : ( n441 ) ;
assign n443 =  ( LB2D_shift_x ) >= ( 9'd8 )  ;
assign n444 =  ( LB2D_shift_x ) == ( 9'd0 )  ;
assign n445 =  ( n443 ) | ( n444 )  ;
assign n446 = n136[71:64] ;
assign n447 = LB2D_shift_7[71:64] ;
assign n448 = LB2D_shift_6[71:64] ;
assign n449 = LB2D_shift_5[71:64] ;
assign n450 = LB2D_shift_4[71:64] ;
assign n451 = LB2D_shift_3[71:64] ;
assign n452 = LB2D_shift_2[71:64] ;
assign n453 = LB2D_shift_1[71:64] ;
assign n454 = LB2D_shift_0[71:64] ;
assign n455 =  { ( n453 ) , ( n454 ) }  ;
assign n456 =  { ( n452 ) , ( n455 ) }  ;
assign n457 =  { ( n451 ) , ( n456 ) }  ;
assign n458 =  { ( n450 ) , ( n457 ) }  ;
assign n459 =  { ( n449 ) , ( n458 ) }  ;
assign n460 =  { ( n448 ) , ( n459 ) }  ;
assign n461 =  { ( n447 ) , ( n460 ) }  ;
assign n462 =  { ( n446 ) , ( n461 ) }  ;
assign n463 = n136[63:56] ;
assign n464 = LB2D_shift_7[63:56] ;
assign n465 = LB2D_shift_6[63:56] ;
assign n466 = LB2D_shift_5[63:56] ;
assign n467 = LB2D_shift_4[63:56] ;
assign n468 = LB2D_shift_3[63:56] ;
assign n469 = LB2D_shift_2[63:56] ;
assign n470 = LB2D_shift_1[63:56] ;
assign n471 = LB2D_shift_0[63:56] ;
assign n472 =  { ( n470 ) , ( n471 ) }  ;
assign n473 =  { ( n469 ) , ( n472 ) }  ;
assign n474 =  { ( n468 ) , ( n473 ) }  ;
assign n475 =  { ( n467 ) , ( n474 ) }  ;
assign n476 =  { ( n466 ) , ( n475 ) }  ;
assign n477 =  { ( n465 ) , ( n476 ) }  ;
assign n478 =  { ( n464 ) , ( n477 ) }  ;
assign n479 =  { ( n463 ) , ( n478 ) }  ;
assign n480 = n136[55:48] ;
assign n481 = LB2D_shift_7[55:48] ;
assign n482 = LB2D_shift_6[55:48] ;
assign n483 = LB2D_shift_5[55:48] ;
assign n484 = LB2D_shift_4[55:48] ;
assign n485 = LB2D_shift_3[55:48] ;
assign n486 = LB2D_shift_2[55:48] ;
assign n487 = LB2D_shift_1[55:48] ;
assign n488 = LB2D_shift_0[55:48] ;
assign n489 =  { ( n487 ) , ( n488 ) }  ;
assign n490 =  { ( n486 ) , ( n489 ) }  ;
assign n491 =  { ( n485 ) , ( n490 ) }  ;
assign n492 =  { ( n484 ) , ( n491 ) }  ;
assign n493 =  { ( n483 ) , ( n492 ) }  ;
assign n494 =  { ( n482 ) , ( n493 ) }  ;
assign n495 =  { ( n481 ) , ( n494 ) }  ;
assign n496 =  { ( n480 ) , ( n495 ) }  ;
assign n497 = n136[47:40] ;
assign n498 = LB2D_shift_7[47:40] ;
assign n499 = LB2D_shift_6[47:40] ;
assign n500 = LB2D_shift_5[47:40] ;
assign n501 = LB2D_shift_4[47:40] ;
assign n502 = LB2D_shift_3[47:40] ;
assign n503 = LB2D_shift_2[47:40] ;
assign n504 = LB2D_shift_1[47:40] ;
assign n505 = LB2D_shift_0[47:40] ;
assign n506 =  { ( n504 ) , ( n505 ) }  ;
assign n507 =  { ( n503 ) , ( n506 ) }  ;
assign n508 =  { ( n502 ) , ( n507 ) }  ;
assign n509 =  { ( n501 ) , ( n508 ) }  ;
assign n510 =  { ( n500 ) , ( n509 ) }  ;
assign n511 =  { ( n499 ) , ( n510 ) }  ;
assign n512 =  { ( n498 ) , ( n511 ) }  ;
assign n513 =  { ( n497 ) , ( n512 ) }  ;
assign n514 = n136[39:32] ;
assign n515 = LB2D_shift_7[39:32] ;
assign n516 = LB2D_shift_6[39:32] ;
assign n517 = LB2D_shift_5[39:32] ;
assign n518 = LB2D_shift_4[39:32] ;
assign n519 = LB2D_shift_3[39:32] ;
assign n520 = LB2D_shift_2[39:32] ;
assign n521 = LB2D_shift_1[39:32] ;
assign n522 = LB2D_shift_0[39:32] ;
assign n523 =  { ( n521 ) , ( n522 ) }  ;
assign n524 =  { ( n520 ) , ( n523 ) }  ;
assign n525 =  { ( n519 ) , ( n524 ) }  ;
assign n526 =  { ( n518 ) , ( n525 ) }  ;
assign n527 =  { ( n517 ) , ( n526 ) }  ;
assign n528 =  { ( n516 ) , ( n527 ) }  ;
assign n529 =  { ( n515 ) , ( n528 ) }  ;
assign n530 =  { ( n514 ) , ( n529 ) }  ;
assign n531 = n136[31:24] ;
assign n532 = LB2D_shift_7[31:24] ;
assign n533 = LB2D_shift_6[31:24] ;
assign n534 = LB2D_shift_5[31:24] ;
assign n535 = LB2D_shift_4[31:24] ;
assign n536 = LB2D_shift_3[31:24] ;
assign n537 = LB2D_shift_2[31:24] ;
assign n538 = LB2D_shift_1[31:24] ;
assign n539 = LB2D_shift_0[31:24] ;
assign n540 =  { ( n538 ) , ( n539 ) }  ;
assign n541 =  { ( n537 ) , ( n540 ) }  ;
assign n542 =  { ( n536 ) , ( n541 ) }  ;
assign n543 =  { ( n535 ) , ( n542 ) }  ;
assign n544 =  { ( n534 ) , ( n543 ) }  ;
assign n545 =  { ( n533 ) , ( n544 ) }  ;
assign n546 =  { ( n532 ) , ( n545 ) }  ;
assign n547 =  { ( n531 ) , ( n546 ) }  ;
assign n548 = n136[23:16] ;
assign n549 = LB2D_shift_7[23:16] ;
assign n550 = LB2D_shift_6[23:16] ;
assign n551 = LB2D_shift_5[23:16] ;
assign n552 = LB2D_shift_4[23:16] ;
assign n553 = LB2D_shift_3[23:16] ;
assign n554 = LB2D_shift_2[23:16] ;
assign n555 = LB2D_shift_1[23:16] ;
assign n556 = LB2D_shift_0[23:16] ;
assign n557 =  { ( n555 ) , ( n556 ) }  ;
assign n558 =  { ( n554 ) , ( n557 ) }  ;
assign n559 =  { ( n553 ) , ( n558 ) }  ;
assign n560 =  { ( n552 ) , ( n559 ) }  ;
assign n561 =  { ( n551 ) , ( n560 ) }  ;
assign n562 =  { ( n550 ) , ( n561 ) }  ;
assign n563 =  { ( n549 ) , ( n562 ) }  ;
assign n564 =  { ( n548 ) , ( n563 ) }  ;
assign n565 = n136[15:8] ;
assign n566 = LB2D_shift_7[15:8] ;
assign n567 = LB2D_shift_6[15:8] ;
assign n568 = LB2D_shift_5[15:8] ;
assign n569 = LB2D_shift_4[15:8] ;
assign n570 = LB2D_shift_3[15:8] ;
assign n571 = LB2D_shift_2[15:8] ;
assign n572 = LB2D_shift_1[15:8] ;
assign n573 = LB2D_shift_0[15:8] ;
assign n574 =  { ( n572 ) , ( n573 ) }  ;
assign n575 =  { ( n571 ) , ( n574 ) }  ;
assign n576 =  { ( n570 ) , ( n575 ) }  ;
assign n577 =  { ( n569 ) , ( n576 ) }  ;
assign n578 =  { ( n568 ) , ( n577 ) }  ;
assign n579 =  { ( n567 ) , ( n578 ) }  ;
assign n580 =  { ( n566 ) , ( n579 ) }  ;
assign n581 =  { ( n565 ) , ( n580 ) }  ;
assign n582 = n136[7:0] ;
assign n583 = LB2D_shift_7[7:0] ;
assign n584 = LB2D_shift_6[7:0] ;
assign n585 = LB2D_shift_5[7:0] ;
assign n586 = LB2D_shift_4[7:0] ;
assign n587 = LB2D_shift_3[7:0] ;
assign n588 = LB2D_shift_2[7:0] ;
assign n589 = LB2D_shift_1[7:0] ;
assign n590 = LB2D_shift_0[7:0] ;
assign n591 =  { ( n589 ) , ( n590 ) }  ;
assign n592 =  { ( n588 ) , ( n591 ) }  ;
assign n593 =  { ( n587 ) , ( n592 ) }  ;
assign n594 =  { ( n586 ) , ( n593 ) }  ;
assign n595 =  { ( n585 ) , ( n594 ) }  ;
assign n596 =  { ( n584 ) , ( n595 ) }  ;
assign n597 =  { ( n583 ) , ( n596 ) }  ;
assign n598 =  { ( n582 ) , ( n597 ) }  ;
assign n599 =  { ( n581 ) , ( n598 ) }  ;
assign n600 =  { ( n564 ) , ( n599 ) }  ;
assign n601 =  { ( n547 ) , ( n600 ) }  ;
assign n602 =  { ( n530 ) , ( n601 ) }  ;
assign n603 =  { ( n513 ) , ( n602 ) }  ;
assign n604 =  { ( n496 ) , ( n603 ) }  ;
assign n605 =  { ( n479 ) , ( n604 ) }  ;
assign n606 =  { ( n462 ) , ( n605 ) }  ;
assign n607 =  ( n445 ) ? ( n606 ) : ( stencil_stream_buff_0 ) ;
assign n608 =  ( n33 ) ? ( stencil_stream_buff_0 ) : ( stencil_stream_buff_0 ) ;
assign n609 =  ( n30 ) ? ( stencil_stream_buff_0 ) : ( n608 ) ;
assign n610 =  ( n25 ) ? ( n607 ) : ( n609 ) ;
assign n611 =  ( n18 ) ? ( stencil_stream_buff_0 ) : ( n610 ) ;
assign n612 =  ( n9 ) ? ( stencil_stream_buff_0 ) : ( n611 ) ;
assign n613 =  ( n4 ) ? ( stencil_stream_buff_0 ) : ( n612 ) ;
assign n614 =  ( n25 ) & ( n445 )  ;
assign n615 =  ( n33 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_1 ) ;
assign n616 =  ( n30 ) ? ( stencil_stream_buff_1 ) : ( n615 ) ;
assign n617 =  ( n614 ) ? ( stencil_stream_buff_0 ) : ( n616 ) ;
assign n618 =  ( n18 ) ? ( stencil_stream_buff_1 ) : ( n617 ) ;
assign n619 =  ( n9 ) ? ( stencil_stream_buff_1 ) : ( n618 ) ;
assign n620 =  ( n4 ) ? ( stencil_stream_buff_1 ) : ( n619 ) ;
assign n621 =  ( n163 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n622 = ~ ( n445 ) ;
assign n623 =  ( n622 ) ? ( stencil_stream_empty ) : ( 1'd0 ) ;
assign n624 =  ( n33 ) ? ( stencil_stream_empty ) : ( stencil_stream_empty ) ;
assign n625 =  ( n30 ) ? ( stencil_stream_empty ) : ( n624 ) ;
assign n626 =  ( n25 ) ? ( n623 ) : ( n625 ) ;
assign n627 =  ( n18 ) ? ( n621 ) : ( n626 ) ;
assign n628 =  ( n9 ) ? ( stencil_stream_empty ) : ( n627 ) ;
assign n629 =  ( n4 ) ? ( stencil_stream_empty ) : ( n628 ) ;
assign n630 =  ( n14 ) ? ( 1'd0 ) : ( 1'd0 ) ;
assign n631 =  ( stencil_stream_empty ) == ( 1'd1 )  ;
assign n632 =  ( n631 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n633 =  ( n622 ) ? ( stencil_stream_full ) : ( n632 ) ;
assign n634 =  ( n33 ) ? ( stencil_stream_full ) : ( stencil_stream_full ) ;
assign n635 =  ( n30 ) ? ( stencil_stream_full ) : ( n634 ) ;
assign n636 =  ( n25 ) ? ( n633 ) : ( n635 ) ;
assign n637 =  ( n18 ) ? ( n630 ) : ( n636 ) ;
assign n638 =  ( n9 ) ? ( stencil_stream_full ) : ( n637 ) ;
assign n639 =  ( n4 ) ? ( stencil_stream_full ) : ( n638 ) ;
assign n640 = ~ ( n4 ) ;
assign n641 =  ( 1'b1 ) & ( n640 )  ;
assign n642 = ~ ( n9 ) ;
assign n643 =  ( n641 ) & ( n642 )  ;
assign n644 = ~ ( n18 ) ;
assign n645 =  ( n643 ) & ( n644 )  ;
assign n646 = ~ ( n25 ) ;
assign n647 =  ( n645 ) & ( n646 )  ;
assign n648 = ~ ( n30 ) ;
assign n649 =  ( n647 ) & ( n648 )  ;
assign n650 = ~ ( n33 ) ;
assign n651 =  ( n649 ) & ( n650 )  ;
assign n652 =  ( n649 ) & ( n33 )  ;
assign n653 =  ( n647 ) & ( n30 )  ;
assign n654 = ~ ( n332 ) ;
assign n655 =  ( n653 ) & ( n654 )  ;
assign n656 =  ( n653 ) & ( n332 )  ;
assign n657 =  ( n645 ) & ( n25 )  ;
assign n658 =  ( n643 ) & ( n18 )  ;
assign n659 =  ( n641 ) & ( n9 )  ;
assign n660 =  ( 1'b1 ) & ( n4 )  ;
assign LB2D_proc_0_addr0 = n656 ? (n333) : (0);
assign LB2D_proc_0_data0 = n656 ? (n331) : ('dx);
assign LB2D_proc_0_wen0 = n656 ? ( 1'b1 ) : (1'b0);
assign n661 = ~ ( n335 ) ;
assign n662 =  ( n653 ) & ( n661 )  ;
assign n663 =  ( n653 ) & ( n335 )  ;
assign LB2D_proc_1_addr0 = n663 ? (n333) : (0);
assign LB2D_proc_1_data0 = n663 ? (n331) : ('dx);
assign LB2D_proc_1_wen0 = n663 ? ( 1'b1 ) : (1'b0);
assign n664 = ~ ( n337 ) ;
assign n665 =  ( n653 ) & ( n664 )  ;
assign n666 =  ( n653 ) & ( n337 )  ;
assign LB2D_proc_2_addr0 = n666 ? (n333) : (0);
assign LB2D_proc_2_data0 = n666 ? (n331) : ('dx);
assign LB2D_proc_2_wen0 = n666 ? ( 1'b1 ) : (1'b0);
assign n667 = ~ ( n339 ) ;
assign n668 =  ( n653 ) & ( n667 )  ;
assign n669 =  ( n653 ) & ( n339 )  ;
assign LB2D_proc_3_addr0 = n669 ? (n333) : (0);
assign LB2D_proc_3_data0 = n669 ? (n331) : ('dx);
assign LB2D_proc_3_wen0 = n669 ? ( 1'b1 ) : (1'b0);
assign n670 = ~ ( n341 ) ;
assign n671 =  ( n653 ) & ( n670 )  ;
assign n672 =  ( n653 ) & ( n341 )  ;
assign LB2D_proc_4_addr0 = n672 ? (n333) : (0);
assign LB2D_proc_4_data0 = n672 ? (n331) : ('dx);
assign LB2D_proc_4_wen0 = n672 ? ( 1'b1 ) : (1'b0);
assign n673 = ~ ( n343 ) ;
assign n674 =  ( n653 ) & ( n673 )  ;
assign n675 =  ( n653 ) & ( n343 )  ;
assign LB2D_proc_5_addr0 = n675 ? (n333) : (0);
assign LB2D_proc_5_data0 = n675 ? (n331) : ('dx);
assign LB2D_proc_5_wen0 = n675 ? ( 1'b1 ) : (1'b0);
assign n676 = ~ ( n345 ) ;
assign n677 =  ( n653 ) & ( n676 )  ;
assign n678 =  ( n653 ) & ( n345 )  ;
assign LB2D_proc_6_addr0 = n678 ? (n333) : (0);
assign LB2D_proc_6_data0 = n678 ? (n331) : ('dx);
assign LB2D_proc_6_wen0 = n678 ? ( 1'b1 ) : (1'b0);
assign n679 = ~ ( n65 ) ;
assign n680 =  ( n653 ) & ( n679 )  ;
assign n681 =  ( n653 ) & ( n65 )  ;
assign LB2D_proc_7_addr0 = n681 ? (n333) : (0);
assign LB2D_proc_7_data0 = n681 ? (n331) : ('dx);
assign LB2D_proc_7_wen0 = n681 ? ( 1'b1 ) : (1'b0);
always @(posedge clk) begin
   if(rst) begin
       LB1D_buff <= LB1D_buff;
       LB1D_in <= LB1D_in;
       LB1D_it_1 <= LB1D_it_1;
       LB1D_p_cnt <= LB1D_p_cnt;
       LB1D_uIn <= LB1D_uIn;
       LB2D_proc_w <= LB2D_proc_w;
       LB2D_proc_x <= LB2D_proc_x;
       LB2D_proc_y <= LB2D_proc_y;
       LB2D_shift_0 <= LB2D_shift_0;
       LB2D_shift_1 <= LB2D_shift_1;
       LB2D_shift_2 <= LB2D_shift_2;
       LB2D_shift_3 <= LB2D_shift_3;
       LB2D_shift_4 <= LB2D_shift_4;
       LB2D_shift_5 <= LB2D_shift_5;
       LB2D_shift_6 <= LB2D_shift_6;
       LB2D_shift_7 <= LB2D_shift_7;
       LB2D_shift_x <= LB2D_shift_x;
       LB2D_shift_y <= LB2D_shift_y;
       arg_0_TDATA <= arg_0_TDATA;
       arg_0_TVALID <= arg_0_TVALID;
       arg_1_TREADY <= arg_1_TREADY;
       gb_exit_it_1 <= gb_exit_it_1;
       gb_exit_it_2 <= gb_exit_it_2;
       gb_exit_it_3 <= gb_exit_it_3;
       gb_exit_it_4 <= gb_exit_it_4;
       gb_exit_it_5 <= gb_exit_it_5;
       gb_exit_it_6 <= gb_exit_it_6;
       gb_exit_it_7 <= gb_exit_it_7;
       gb_exit_it_8 <= gb_exit_it_8;
       gb_p_cnt <= gb_p_cnt;
       gb_pp_it_1 <= gb_pp_it_1;
       gb_pp_it_2 <= gb_pp_it_2;
       gb_pp_it_3 <= gb_pp_it_3;
       gb_pp_it_4 <= gb_pp_it_4;
       gb_pp_it_5 <= gb_pp_it_5;
       gb_pp_it_6 <= gb_pp_it_6;
       gb_pp_it_7 <= gb_pp_it_7;
       gb_pp_it_8 <= gb_pp_it_8;
       gb_pp_it_9 <= gb_pp_it_9;
       in_stream_buff_0 <= in_stream_buff_0;
       in_stream_buff_1 <= in_stream_buff_1;
       in_stream_empty <= in_stream_empty;
       in_stream_full <= in_stream_full;
       slice_stream_buff_0 <= slice_stream_buff_0;
       slice_stream_buff_1 <= slice_stream_buff_1;
       slice_stream_empty <= slice_stream_empty;
       slice_stream_full <= slice_stream_full;
       stencil_stream_buff_0 <= stencil_stream_buff_0;
       stencil_stream_buff_1 <= stencil_stream_buff_1;
       stencil_stream_empty <= stencil_stream_empty;
       stencil_stream_full <= stencil_stream_full;
   end
   else if(step) begin
       LB1D_buff <= n39;
       LB1D_in <= n45;
       LB1D_it_1 <= n50;
       LB1D_p_cnt <= n58;
       LB1D_uIn <= n63;
       LB2D_proc_w <= n74;
       LB2D_proc_x <= n82;
       LB2D_proc_y <= n92;
       LB2D_shift_0 <= n98;
       LB2D_shift_1 <= n104;
       LB2D_shift_2 <= n110;
       LB2D_shift_3 <= n116;
       LB2D_shift_4 <= n122;
       LB2D_shift_5 <= n128;
       LB2D_shift_6 <= n134;
       LB2D_shift_7 <= n142;
       LB2D_shift_x <= n151;
       LB2D_shift_y <= n162;
       arg_0_TDATA <= n173;
       arg_0_TVALID <= n183;
       arg_1_TREADY <= n189;
       gb_exit_it_1 <= n197;
       gb_exit_it_2 <= n203;
       gb_exit_it_3 <= n209;
       gb_exit_it_4 <= n215;
       gb_exit_it_5 <= n221;
       gb_exit_it_6 <= n227;
       gb_exit_it_7 <= n233;
       gb_exit_it_8 <= n239;
       gb_p_cnt <= n248;
       gb_pp_it_1 <= n254;
       gb_pp_it_2 <= n260;
       gb_pp_it_3 <= n266;
       gb_pp_it_4 <= n272;
       gb_pp_it_5 <= n278;
       gb_pp_it_6 <= n284;
       gb_pp_it_7 <= n290;
       gb_pp_it_8 <= n296;
       gb_pp_it_9 <= n302;
       in_stream_buff_0 <= n308;
       in_stream_buff_1 <= n314;
       in_stream_empty <= n322;
       in_stream_full <= n330;
       slice_stream_buff_0 <= n418;
       slice_stream_buff_1 <= n425;
       slice_stream_empty <= n433;
       slice_stream_full <= n442;
       stencil_stream_buff_0 <= n613;
       stencil_stream_buff_1 <= n620;
       stencil_stream_empty <= n629;
       stencil_stream_full <= n639;
       if (LB2D_proc_0_wen0) begin
           LB2D_proc_0 [ LB2D_proc_0_addr0 ] <= LB2D_proc_0_data0 ;
       end
       if (LB2D_proc_1_wen0) begin
           LB2D_proc_1 [ LB2D_proc_1_addr0 ] <= LB2D_proc_1_data0 ;
       end
       if (LB2D_proc_2_wen0) begin
           LB2D_proc_2 [ LB2D_proc_2_addr0 ] <= LB2D_proc_2_data0 ;
       end
       if (LB2D_proc_3_wen0) begin
           LB2D_proc_3 [ LB2D_proc_3_addr0 ] <= LB2D_proc_3_data0 ;
       end
       if (LB2D_proc_4_wen0) begin
           LB2D_proc_4 [ LB2D_proc_4_addr0 ] <= LB2D_proc_4_data0 ;
       end
       if (LB2D_proc_5_wen0) begin
           LB2D_proc_5 [ LB2D_proc_5_addr0 ] <= LB2D_proc_5_data0 ;
       end
       if (LB2D_proc_6_wen0) begin
           LB2D_proc_6 [ LB2D_proc_6_addr0 ] <= LB2D_proc_6_data0 ;
       end
       if (LB2D_proc_7_wen0) begin
           LB2D_proc_7 [ LB2D_proc_7_addr0 ] <= LB2D_proc_7_data0 ;
       end
   end
end
endmodule
