module GB(
arg_0_TREADY,
arg_1_TDATA,
arg_1_TVALID,
LB1D_buff,
LB1D_in,
LB1D_it_1,
LB1D_p_cnt,
LB2D_proc_w,
LB2D_proc_x,
LB2D_proc_y,
LB2D_shift_0,
LB2D_shift_1,
LB2D_shift_2,
LB2D_shift_3,
LB2D_shift_4,
LB2D_shift_5,
LB2D_shift_6,
LB2D_shift_7,
LB2D_shift_x,
LB2D_shift_y,
arg_0_TDATA,
arg_0_TVALID,
arg_1_TREADY,
gb_exit_it_1,
gb_exit_it_2,
gb_exit_it_3,
gb_exit_it_4,
gb_exit_it_5,
gb_exit_it_6,
gb_exit_it_7,
gb_exit_it_8,
gb_p_cnt,
gb_pp_it_1,
gb_pp_it_2,
gb_pp_it_3,
gb_pp_it_4,
gb_pp_it_5,
gb_pp_it_6,
gb_pp_it_7,
gb_pp_it_8,
gb_pp_it_9,
in_stream_buff_0,
in_stream_buff_1,
in_stream_empty,
in_stream_full,
slice_stream_buff_0,
slice_stream_buff_1,
slice_stream_empty,
slice_stream_full,
stencil_stream_buff_0,
stencil_stream_buff_1,
stencil_stream_empty,
stencil_stream_full,
clk,rst,
step
);
input            arg_0_TREADY;
input      [7:0] arg_1_TDATA;
input            arg_1_TVALID;
input clk;
input rst;
input step;
output      [7:0] LB1D_buff;
output      [7:0] LB1D_in;
output            LB1D_it_1;
output     [18:0] LB1D_p_cnt;
output     [63:0] LB2D_proc_w;
output      [8:0] LB2D_proc_x;
output      [9:0] LB2D_proc_y;
output     [71:0] LB2D_shift_0;
output     [71:0] LB2D_shift_1;
output     [71:0] LB2D_shift_2;
output     [71:0] LB2D_shift_3;
output     [71:0] LB2D_shift_4;
output     [71:0] LB2D_shift_5;
output     [71:0] LB2D_shift_6;
output     [71:0] LB2D_shift_7;
output      [8:0] LB2D_shift_x;
output      [9:0] LB2D_shift_y;
output      [7:0] arg_0_TDATA;
output            arg_0_TVALID;
output            arg_1_TREADY;
output            gb_exit_it_1;
output            gb_exit_it_2;
output            gb_exit_it_3;
output            gb_exit_it_4;
output            gb_exit_it_5;
output            gb_exit_it_6;
output            gb_exit_it_7;
output            gb_exit_it_8;
output     [18:0] gb_p_cnt;
output            gb_pp_it_1;
output            gb_pp_it_2;
output            gb_pp_it_3;
output            gb_pp_it_4;
output            gb_pp_it_5;
output            gb_pp_it_6;
output            gb_pp_it_7;
output            gb_pp_it_8;
output            gb_pp_it_9;
output      [7:0] in_stream_buff_0;
output      [7:0] in_stream_buff_1;
output            in_stream_empty;
output            in_stream_full;
output     [71:0] slice_stream_buff_0;
output     [71:0] slice_stream_buff_1;
output            slice_stream_empty;
output            slice_stream_full;
output    [647:0] stencil_stream_buff_0;
output    [647:0] stencil_stream_buff_1;
output            stencil_stream_empty;
output            stencil_stream_full;
reg      [7:0] LB1D_buff;
reg      [7:0] LB1D_in;
reg            LB1D_it_1;
reg     [18:0] LB1D_p_cnt;
reg     [63:0] LB2D_proc_w;
reg      [8:0] LB2D_proc_x;
reg      [9:0] LB2D_proc_y;
reg     [71:0] LB2D_shift_0;
reg     [71:0] LB2D_shift_1;
reg     [71:0] LB2D_shift_2;
reg     [71:0] LB2D_shift_3;
reg     [71:0] LB2D_shift_4;
reg     [71:0] LB2D_shift_5;
reg     [71:0] LB2D_shift_6;
reg     [71:0] LB2D_shift_7;
reg      [8:0] LB2D_shift_x;
reg      [9:0] LB2D_shift_y;
reg      [7:0] arg_0_TDATA;
reg            arg_0_TVALID;
reg            arg_1_TREADY;
reg            gb_exit_it_1;
reg            gb_exit_it_2;
reg            gb_exit_it_3;
reg            gb_exit_it_4;
reg            gb_exit_it_5;
reg            gb_exit_it_6;
reg            gb_exit_it_7;
reg            gb_exit_it_8;
reg     [18:0] gb_p_cnt;
reg            gb_pp_it_1;
reg            gb_pp_it_2;
reg            gb_pp_it_3;
reg            gb_pp_it_4;
reg            gb_pp_it_5;
reg            gb_pp_it_6;
reg            gb_pp_it_7;
reg            gb_pp_it_8;
reg            gb_pp_it_9;
reg      [7:0] in_stream_buff_0;
reg      [7:0] in_stream_buff_1;
reg            in_stream_empty;
reg            in_stream_full;
reg     [71:0] slice_stream_buff_0;
reg     [71:0] slice_stream_buff_1;
reg            slice_stream_empty;
reg            slice_stream_full;
reg    [647:0] stencil_stream_buff_0;
reg    [647:0] stencil_stream_buff_1;
reg            stencil_stream_empty;
reg            stencil_stream_full;
wire            arg_0_TREADY;
wire      [7:0] arg_1_TDATA;
wire            arg_1_TVALID;
wire            n0;
wire            n1;
wire            n2;
wire            n3;
wire            n4;
wire            n5;
wire            n6;
wire            n7;
wire            n8;
wire            n9;
wire            n10;
wire            n11;
wire            n12;
wire            n13;
wire            n14;
wire            n15;
wire            n16;
wire            n17;
wire            n18;
wire            n19;
wire            n20;
wire            n21;
wire            n22;
wire            n23;
wire            n24;
wire            n25;
wire            n26;
wire            n27;
wire            n28;
wire            n29;
wire            n30;
wire            n31;
wire            n32;
wire            n33;
wire            n34;
wire            n35;
wire            n36;
wire            n37;
wire      [7:0] n38;
wire      [7:0] n39;
wire      [7:0] n40;
wire      [7:0] n41;
wire      [7:0] n42;
wire      [7:0] n43;
wire      [7:0] n44;
wire      [7:0] n45;
wire            n46;
wire            n47;
wire            n48;
wire     [18:0] n49;
wire     [18:0] n50;
wire            n51;
wire     [18:0] n52;
wire     [18:0] n53;
wire     [18:0] n54;
wire     [18:0] n55;
wire     [18:0] n56;
wire     [18:0] n57;
wire     [18:0] n58;
wire     [18:0] n59;
wire            n60;
wire            n61;
wire     [63:0] n62;
wire     [63:0] n63;
wire     [63:0] n64;
wire     [63:0] n65;
wire     [63:0] n66;
wire     [63:0] n67;
wire     [63:0] n68;
wire     [63:0] n69;
wire     [63:0] n70;
wire            n71;
wire            n72;
wire            n73;
wire      [8:0] n74;
wire      [8:0] n75;
wire      [8:0] n76;
wire      [8:0] n77;
wire      [8:0] n78;
wire      [8:0] n79;
wire      [8:0] n80;
wire      [8:0] n81;
wire            n82;
wire      [9:0] n83;
wire      [9:0] n84;
wire      [9:0] n85;
wire      [9:0] n86;
wire      [9:0] n87;
wire      [9:0] n88;
wire      [9:0] n89;
wire            n90;
wire     [71:0] n91;
wire     [71:0] n92;
wire     [71:0] n93;
wire     [71:0] n94;
wire     [71:0] n95;
wire     [71:0] n96;
wire     [71:0] n97;
wire     [71:0] n98;
wire     [71:0] n99;
wire     [71:0] n100;
wire     [71:0] n101;
wire     [71:0] n102;
wire     [71:0] n103;
wire     [71:0] n104;
wire     [71:0] n105;
wire     [71:0] n106;
wire     [71:0] n107;
wire     [71:0] n108;
wire     [71:0] n109;
wire     [71:0] n110;
wire     [71:0] n111;
wire     [71:0] n112;
wire     [71:0] n113;
wire     [71:0] n114;
wire     [71:0] n115;
wire     [71:0] n116;
wire     [71:0] n117;
wire     [71:0] n118;
wire     [71:0] n119;
wire     [71:0] n120;
wire     [71:0] n121;
wire     [71:0] n122;
wire     [71:0] n123;
wire     [71:0] n124;
wire     [71:0] n125;
wire     [71:0] n126;
wire     [71:0] n127;
wire     [71:0] n128;
wire     [71:0] n129;
wire     [71:0] n130;
wire     [71:0] n131;
wire     [71:0] n132;
wire     [71:0] n133;
wire     [71:0] n134;
wire     [71:0] n135;
wire     [71:0] n136;
wire     [71:0] n137;
wire     [71:0] n138;
wire     [71:0] n139;
wire      [8:0] n140;
wire      [8:0] n141;
wire      [8:0] n142;
wire      [8:0] n143;
wire      [8:0] n144;
wire      [8:0] n145;
wire      [8:0] n146;
wire            n147;
wire            n148;
wire      [9:0] n149;
wire      [9:0] n150;
wire      [9:0] n151;
wire      [9:0] n152;
wire      [9:0] n153;
wire      [9:0] n154;
wire      [9:0] n155;
wire      [9:0] n156;
wire      [9:0] n157;
wire            n158;
wire    [647:0] n159;
wire      [7:0] n160;
wire      [7:0] n161;
wire      [7:0] n162;
wire      [7:0] n163;
wire      [7:0] n164;
wire      [7:0] n165;
wire      [7:0] n166;
wire            n167;
wire            n168;
wire            n169;
wire            n170;
wire            n171;
wire            n172;
wire            n173;
wire            n174;
wire            n175;
wire            n176;
wire            n177;
wire            n178;
wire            n179;
wire            n180;
wire            n181;
wire     [18:0] n182;
wire            n183;
wire            n184;
wire            n185;
wire            n186;
wire            n187;
wire            n188;
wire            n189;
wire            n190;
wire            n191;
wire            n192;
wire            n193;
wire            n194;
wire            n195;
wire            n196;
wire            n197;
wire            n198;
wire            n199;
wire            n200;
wire            n201;
wire            n202;
wire            n203;
wire            n204;
wire            n205;
wire            n206;
wire            n207;
wire            n208;
wire            n209;
wire            n210;
wire            n211;
wire            n212;
wire            n213;
wire            n214;
wire            n215;
wire            n216;
wire            n217;
wire            n218;
wire            n219;
wire            n220;
wire            n221;
wire            n222;
wire            n223;
wire            n224;
wire            n225;
wire            n226;
wire            n227;
wire            n228;
wire            n229;
wire            n230;
wire            n231;
wire            n232;
wire            n233;
wire     [18:0] n234;
wire     [18:0] n235;
wire     [18:0] n236;
wire     [18:0] n237;
wire     [18:0] n238;
wire     [18:0] n239;
wire     [18:0] n240;
wire            n241;
wire            n242;
wire            n243;
wire            n244;
wire            n245;
wire            n246;
wire            n247;
wire            n248;
wire            n249;
wire            n250;
wire            n251;
wire            n252;
wire            n253;
wire            n254;
wire            n255;
wire            n256;
wire            n257;
wire            n258;
wire            n259;
wire            n260;
wire            n261;
wire            n262;
wire            n263;
wire            n264;
wire            n265;
wire            n266;
wire            n267;
wire            n268;
wire            n269;
wire            n270;
wire            n271;
wire            n272;
wire            n273;
wire            n274;
wire            n275;
wire            n276;
wire            n277;
wire            n278;
wire            n279;
wire            n280;
wire            n281;
wire            n282;
wire            n283;
wire            n284;
wire            n285;
wire            n286;
wire            n287;
wire            n288;
wire            n289;
wire            n290;
wire            n291;
wire            n292;
wire            n293;
wire            n294;
wire      [7:0] n295;
wire      [7:0] n296;
wire      [7:0] n297;
wire      [7:0] n298;
wire      [7:0] n299;
wire      [7:0] n300;
wire      [7:0] n301;
wire      [7:0] n302;
wire      [7:0] n303;
wire      [7:0] n304;
wire      [7:0] n305;
wire      [7:0] n306;
wire            n307;
wire            n308;
wire            n309;
wire            n310;
wire            n311;
wire            n312;
wire            n313;
wire            n314;
wire            n315;
wire            n316;
wire            n317;
wire            n318;
wire            n319;
wire            n320;
wire            n321;
wire            n322;
wire      [7:0] n323;
wire            n324;
wire      [7:0] n325;
wire            n326;
wire      [7:0] n327;
wire            n328;
wire      [7:0] n329;
wire            n330;
wire      [7:0] n331;
wire            n332;
wire      [7:0] n333;
wire            n334;
wire      [7:0] n335;
wire            n336;
wire      [7:0] n337;
wire      [7:0] n338;
wire      [7:0] n339;
wire      [7:0] n340;
wire      [7:0] n341;
wire      [7:0] n342;
wire      [7:0] n343;
wire      [7:0] n344;
wire      [7:0] n345;
wire      [7:0] n346;
wire      [7:0] n347;
wire      [7:0] n348;
wire      [7:0] n349;
wire      [7:0] n350;
wire      [7:0] n351;
wire      [7:0] n352;
wire      [7:0] n353;
wire      [7:0] n354;
wire      [7:0] n355;
wire      [7:0] n356;
wire      [7:0] n357;
wire      [7:0] n358;
wire      [7:0] n359;
wire      [7:0] n360;
wire      [7:0] n361;
wire      [7:0] n362;
wire      [7:0] n363;
wire      [7:0] n364;
wire      [7:0] n365;
wire      [7:0] n366;
wire      [7:0] n367;
wire      [7:0] n368;
wire      [7:0] n369;
wire      [7:0] n370;
wire      [7:0] n371;
wire      [7:0] n372;
wire      [7:0] n373;
wire      [7:0] n374;
wire      [7:0] n375;
wire      [7:0] n376;
wire      [7:0] n377;
wire      [7:0] n378;
wire      [7:0] n379;
wire      [7:0] n380;
wire      [7:0] n381;
wire      [7:0] n382;
wire      [7:0] n383;
wire      [7:0] n384;
wire      [7:0] n385;
wire      [7:0] n386;
wire      [7:0] n387;
wire      [7:0] n388;
wire      [7:0] n389;
wire      [7:0] n390;
wire      [7:0] n391;
wire      [7:0] n392;
wire      [7:0] n393;
wire      [7:0] n394;
wire     [15:0] n395;
wire     [23:0] n396;
wire     [31:0] n397;
wire     [39:0] n398;
wire     [47:0] n399;
wire     [55:0] n400;
wire     [63:0] n401;
wire     [71:0] n402;
wire     [71:0] n403;
wire     [71:0] n404;
wire     [71:0] n405;
wire     [71:0] n406;
wire     [71:0] n407;
wire     [71:0] n408;
wire     [71:0] n409;
wire     [71:0] n410;
wire     [71:0] n411;
wire     [71:0] n412;
wire     [71:0] n413;
wire     [71:0] n414;
wire     [71:0] n415;
wire     [71:0] n416;
wire            n417;
wire            n418;
wire            n419;
wire            n420;
wire            n421;
wire            n422;
wire            n423;
wire            n424;
wire            n425;
wire            n426;
wire            n427;
wire            n428;
wire            n429;
wire            n430;
wire            n431;
wire            n432;
wire            n433;
wire            n434;
wire      [7:0] n435;
wire      [7:0] n436;
wire      [7:0] n437;
wire      [7:0] n438;
wire      [7:0] n439;
wire      [7:0] n440;
wire      [7:0] n441;
wire      [7:0] n442;
wire      [7:0] n443;
wire     [15:0] n444;
wire     [23:0] n445;
wire     [31:0] n446;
wire     [39:0] n447;
wire     [47:0] n448;
wire     [55:0] n449;
wire     [63:0] n450;
wire     [71:0] n451;
wire      [7:0] n452;
wire      [7:0] n453;
wire      [7:0] n454;
wire      [7:0] n455;
wire      [7:0] n456;
wire      [7:0] n457;
wire      [7:0] n458;
wire      [7:0] n459;
wire      [7:0] n460;
wire     [15:0] n461;
wire     [23:0] n462;
wire     [31:0] n463;
wire     [39:0] n464;
wire     [47:0] n465;
wire     [55:0] n466;
wire     [63:0] n467;
wire     [71:0] n468;
wire      [7:0] n469;
wire      [7:0] n470;
wire      [7:0] n471;
wire      [7:0] n472;
wire      [7:0] n473;
wire      [7:0] n474;
wire      [7:0] n475;
wire      [7:0] n476;
wire      [7:0] n477;
wire     [15:0] n478;
wire     [23:0] n479;
wire     [31:0] n480;
wire     [39:0] n481;
wire     [47:0] n482;
wire     [55:0] n483;
wire     [63:0] n484;
wire     [71:0] n485;
wire      [7:0] n486;
wire      [7:0] n487;
wire      [7:0] n488;
wire      [7:0] n489;
wire      [7:0] n490;
wire      [7:0] n491;
wire      [7:0] n492;
wire      [7:0] n493;
wire      [7:0] n494;
wire     [15:0] n495;
wire     [23:0] n496;
wire     [31:0] n497;
wire     [39:0] n498;
wire     [47:0] n499;
wire     [55:0] n500;
wire     [63:0] n501;
wire     [71:0] n502;
wire      [7:0] n503;
wire      [7:0] n504;
wire      [7:0] n505;
wire      [7:0] n506;
wire      [7:0] n507;
wire      [7:0] n508;
wire      [7:0] n509;
wire      [7:0] n510;
wire      [7:0] n511;
wire     [15:0] n512;
wire     [23:0] n513;
wire     [31:0] n514;
wire     [39:0] n515;
wire     [47:0] n516;
wire     [55:0] n517;
wire     [63:0] n518;
wire     [71:0] n519;
wire      [7:0] n520;
wire      [7:0] n521;
wire      [7:0] n522;
wire      [7:0] n523;
wire      [7:0] n524;
wire      [7:0] n525;
wire      [7:0] n526;
wire      [7:0] n527;
wire      [7:0] n528;
wire     [15:0] n529;
wire     [23:0] n530;
wire     [31:0] n531;
wire     [39:0] n532;
wire     [47:0] n533;
wire     [55:0] n534;
wire     [63:0] n535;
wire     [71:0] n536;
wire      [7:0] n537;
wire      [7:0] n538;
wire      [7:0] n539;
wire      [7:0] n540;
wire      [7:0] n541;
wire      [7:0] n542;
wire      [7:0] n543;
wire      [7:0] n544;
wire      [7:0] n545;
wire     [15:0] n546;
wire     [23:0] n547;
wire     [31:0] n548;
wire     [39:0] n549;
wire     [47:0] n550;
wire     [55:0] n551;
wire     [63:0] n552;
wire     [71:0] n553;
wire      [7:0] n554;
wire      [7:0] n555;
wire      [7:0] n556;
wire      [7:0] n557;
wire      [7:0] n558;
wire      [7:0] n559;
wire      [7:0] n560;
wire      [7:0] n561;
wire      [7:0] n562;
wire     [15:0] n563;
wire     [23:0] n564;
wire     [31:0] n565;
wire     [39:0] n566;
wire     [47:0] n567;
wire     [55:0] n568;
wire     [63:0] n569;
wire     [71:0] n570;
wire      [7:0] n571;
wire      [7:0] n572;
wire      [7:0] n573;
wire      [7:0] n574;
wire      [7:0] n575;
wire      [7:0] n576;
wire      [7:0] n577;
wire      [7:0] n578;
wire      [7:0] n579;
wire     [15:0] n580;
wire     [23:0] n581;
wire     [31:0] n582;
wire     [39:0] n583;
wire     [47:0] n584;
wire     [55:0] n585;
wire     [63:0] n586;
wire     [71:0] n587;
wire    [143:0] n588;
wire    [215:0] n589;
wire    [287:0] n590;
wire    [359:0] n591;
wire    [431:0] n592;
wire    [503:0] n593;
wire    [575:0] n594;
wire    [647:0] n595;
wire    [647:0] n596;
wire    [647:0] n597;
wire    [647:0] n598;
wire    [647:0] n599;
wire    [647:0] n600;
wire    [647:0] n601;
wire    [647:0] n602;
wire    [647:0] n603;
wire    [647:0] n604;
wire    [647:0] n605;
wire    [647:0] n606;
wire    [647:0] n607;
wire    [647:0] n608;
wire            n609;
wire            n610;
wire            n611;
wire            n612;
wire            n613;
wire            n614;
wire            n615;
wire            n616;
wire            n617;
wire            n618;
wire            n619;
wire            n620;
wire            n621;
wire            n622;
wire            n623;
wire            n624;
wire            n625;
wire            n626;
wire      [8:0] LB2D_proc_0_addr0;
wire      [7:0] LB2D_proc_0_data0;
wire            n627;
wire            n628;
wire            n629;
wire            n630;
wire            n631;
wire            n632;
wire            n633;
wire            n634;
wire            n635;
wire            n636;
wire            n637;
wire            n638;
wire            n639;
wire            n640;
wire            n641;
wire            n642;
wire            n643;
wire            n644;
wire            n645;
wire      [8:0] LB2D_proc_1_addr0;
wire      [7:0] LB2D_proc_1_data0;
wire            n646;
wire            n647;
wire            n648;
wire      [8:0] LB2D_proc_2_addr0;
wire      [7:0] LB2D_proc_2_data0;
wire            n649;
wire            n650;
wire            n651;
wire      [8:0] LB2D_proc_3_addr0;
wire      [7:0] LB2D_proc_3_data0;
wire            n652;
wire            n653;
wire            n654;
wire      [8:0] LB2D_proc_4_addr0;
wire      [7:0] LB2D_proc_4_data0;
wire            n655;
wire            n656;
wire            n657;
wire      [8:0] LB2D_proc_5_addr0;
wire      [7:0] LB2D_proc_5_data0;
wire            n658;
wire            n659;
wire            n660;
wire      [8:0] LB2D_proc_6_addr0;
wire      [7:0] LB2D_proc_6_data0;
wire            n661;
wire            n662;
wire            n663;
wire      [8:0] LB2D_proc_7_addr0;
wire      [7:0] LB2D_proc_7_data0;
wire            n664;
wire            n665;
wire            n666;
wire            n667;
reg      [7:0] LB2D_proc_0[511:0];
reg      [7:0] LB2D_proc_1[511:0];
reg      [7:0] LB2D_proc_2[511:0];
reg      [7:0] LB2D_proc_3[511:0];
reg      [7:0] LB2D_proc_4[511:0];
reg      [7:0] LB2D_proc_5[511:0];
reg      [7:0] LB2D_proc_6[511:0];
reg      [7:0] LB2D_proc_7[511:0];
wire clk;
wire rst;
wire step;
assign n0 =  ( arg_0_TREADY ) == ( 1'd1 )  ;
assign n1 =  ( arg_0_TVALID ) == ( 1'd1 )  ;
assign n2 =  ( n0 ) & ( n1 )  ;
assign n3 =  ( arg_1_TVALID ) == ( 1'd0 )  ;
assign n4 =  ( n2 ) & ( n3 )  ;
assign n5 =  ( arg_1_TREADY ) == ( 1'd1 )  ;
assign n6 =  ( arg_1_TVALID ) == ( 1'd1 )  ;
assign n7 =  ( n5 ) & ( n6 )  ;
assign n8 =  ( arg_0_TREADY ) == ( 1'd0 )  ;
assign n9 =  ( n7 ) & ( n8 )  ;
assign n10 =  ( arg_0_TVALID ) == ( 1'd0 )  ;
assign n11 =  ( gb_exit_it_1 ) == ( 1'd0 )  ;
assign n12 =  ( stencil_stream_empty ) == ( 1'd0 )  ;
assign n13 =  ( n11 ) & ( n12 )  ;
assign n14 =  ( gb_exit_it_1 ) == ( 1'd1 )  ;
assign n15 =  ( gb_exit_it_8 ) == ( 1'd0 )  ;
assign n16 =  ( n14 ) & ( n15 )  ;
assign n17 =  ( n13 ) | ( n16 )  ;
assign n18 =  ( n10 ) & ( n17 )  ;
assign n19 =  ( slice_stream_empty ) == ( 1'd0 )  ;
assign n20 =  ( LB2D_shift_x ) != ( 9'd488 )  ;
assign n21 =  ( n19 ) & ( n20 )  ;
assign n22 =  ( stencil_stream_full ) == ( 1'd0 )  ;
assign n23 =  ( LB2D_shift_x ) < ( 9'd8 )  ;
assign n24 =  ( n22 ) | ( n23 )  ;
assign n25 =  ( n21 ) & ( n24 )  ;
assign n26 =  ( in_stream_empty ) == ( 1'd0 )  ;
assign n27 =  ( LB2D_proc_x ) != ( 9'd488 )  ;
assign n28 =  ( n26 ) & ( n27 )  ;
assign n29 =  ( slice_stream_full ) == ( 1'd0 )  ;
assign n30 =  ( LB2D_proc_y ) < ( 10'd8 )  ;
assign n31 =  ( n29 ) | ( n30 )  ;
assign n32 =  ( n28 ) & ( n31 )  ;
assign n33 =  ( arg_1_TREADY ) == ( 1'd0 )  ;
assign n34 =  ( in_stream_full ) == ( 1'd0 )  ;
assign n35 =  ( n33 ) & ( n34 )  ;
assign n36 =  ( LB1D_it_1 ) == ( 1'd1 )  ;
assign n37 =  ( n35 ) & ( n36 )  ;
assign n38 =  ( n37 ) ? ( LB1D_in ) : ( LB1D_buff ) ;
assign n39 =  ( n32 ) ? ( LB1D_buff ) : ( n38 ) ;
assign n40 =  ( n25 ) ? ( LB1D_buff ) : ( n39 ) ;
assign n41 =  ( n18 ) ? ( LB1D_buff ) : ( n40 ) ;
assign n42 =  ( n9 ) ? ( LB1D_buff ) : ( n41 ) ;
assign n43 =  ( n4 ) ? ( arg_1_TDATA ) : ( n42 ) ;
assign n44 =  ( n37 ) ? ( LB1D_in ) : ( LB1D_in ) ;
assign n45 =  ( n9 ) ? ( arg_1_TDATA ) : ( n44 ) ;
assign n46 =  ( LB1D_it_1 ) == ( 1'd0 )  ;
assign n47 =  ( n35 ) & ( n46 )  ;
assign n48 =  ( n47 ) ? ( 1'd1 ) : ( LB1D_it_1 ) ;
assign n49 =  ( LB1D_p_cnt ) + ( 19'd1 )  ;
assign n50 =  ( 19'd316224 ) - ( 19'd1 )  ;
assign n51 =  ( LB1D_p_cnt ) == ( n50 )  ;
assign n52 =  ( n51 ) ? ( 19'd0 ) : ( n49 ) ;
assign n53 =  ( n37 ) ? ( n52 ) : ( LB1D_p_cnt ) ;
assign n54 =  ( n47 ) ? ( n49 ) : ( n53 ) ;
assign n55 =  ( n32 ) ? ( LB1D_p_cnt ) : ( n54 ) ;
assign n56 =  ( n25 ) ? ( LB1D_p_cnt ) : ( n55 ) ;
assign n57 =  ( n18 ) ? ( LB1D_p_cnt ) : ( n56 ) ;
assign n58 =  ( n9 ) ? ( LB1D_p_cnt ) : ( n57 ) ;
assign n59 =  ( n4 ) ? ( LB1D_p_cnt ) : ( n58 ) ;
assign n60 =  ( LB2D_proc_w ) < ( 64'd7 )  ;
assign n61 =  ( LB2D_proc_x ) < ( 9'd488 )  ;
assign n62 =  ( LB2D_proc_w ) + ( 64'd1 )  ;
assign n63 =  ( n61 ) ? ( LB2D_proc_w ) : ( n62 ) ;
assign n64 =  ( n60 ) ? ( n63 ) : ( 64'd0 ) ;
assign n65 =  ( n37 ) ? ( LB2D_proc_w ) : ( LB2D_proc_w ) ;
assign n66 =  ( n32 ) ? ( n64 ) : ( n65 ) ;
assign n67 =  ( n25 ) ? ( LB2D_proc_w ) : ( n66 ) ;
assign n68 =  ( n18 ) ? ( LB2D_proc_w ) : ( n67 ) ;
assign n69 =  ( n9 ) ? ( LB2D_proc_w ) : ( n68 ) ;
assign n70 =  ( n4 ) ? ( LB2D_proc_w ) : ( n69 ) ;
assign n71 =  ( LB2D_proc_x ) == ( 9'd488 )  ;
assign n72 =  ( n26 ) & ( n71 )  ;
assign n73 =  ( n72 ) & ( n31 )  ;
assign n74 =  ( LB2D_proc_x ) + ( 9'd1 )  ;
assign n75 =  ( n37 ) ? ( LB2D_proc_x ) : ( LB2D_proc_x ) ;
assign n76 =  ( n32 ) ? ( n74 ) : ( n75 ) ;
assign n77 =  ( n73 ) ? ( 9'd0 ) : ( n76 ) ;
assign n78 =  ( n25 ) ? ( LB2D_proc_x ) : ( n77 ) ;
assign n79 =  ( n18 ) ? ( LB2D_proc_x ) : ( n78 ) ;
assign n80 =  ( n9 ) ? ( LB2D_proc_x ) : ( n79 ) ;
assign n81 =  ( n4 ) ? ( LB2D_proc_x ) : ( n80 ) ;
assign n82 =  ( LB2D_proc_y ) < ( 10'd488 )  ;
assign n83 =  ( n82 ) ? ( LB2D_proc_y ) : ( 10'd488 ) ;
assign n84 =  ( n37 ) ? ( LB2D_proc_y ) : ( LB2D_proc_y ) ;
assign n85 =  ( n32 ) ? ( n83 ) : ( n84 ) ;
assign n86 =  ( n25 ) ? ( LB2D_proc_y ) : ( n85 ) ;
assign n87 =  ( n18 ) ? ( LB2D_proc_y ) : ( n86 ) ;
assign n88 =  ( n9 ) ? ( LB2D_proc_y ) : ( n87 ) ;
assign n89 =  ( n4 ) ? ( LB2D_proc_y ) : ( n88 ) ;
assign n90 =  ( slice_stream_full ) == ( 1'd1 )  ;
assign n91 =  ( n90 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n92 =  ( n37 ) ? ( LB2D_shift_0 ) : ( LB2D_shift_0 ) ;
assign n93 =  ( n32 ) ? ( LB2D_shift_0 ) : ( n92 ) ;
assign n94 =  ( n25 ) ? ( n91 ) : ( n93 ) ;
assign n95 =  ( n18 ) ? ( LB2D_shift_0 ) : ( n94 ) ;
assign n96 =  ( n9 ) ? ( LB2D_shift_0 ) : ( n95 ) ;
assign n97 =  ( n4 ) ? ( LB2D_shift_0 ) : ( n96 ) ;
assign n98 =  ( n37 ) ? ( LB2D_shift_1 ) : ( LB2D_shift_1 ) ;
assign n99 =  ( n32 ) ? ( LB2D_shift_1 ) : ( n98 ) ;
assign n100 =  ( n25 ) ? ( LB2D_shift_0 ) : ( n99 ) ;
assign n101 =  ( n18 ) ? ( LB2D_shift_1 ) : ( n100 ) ;
assign n102 =  ( n9 ) ? ( LB2D_shift_1 ) : ( n101 ) ;
assign n103 =  ( n4 ) ? ( LB2D_shift_1 ) : ( n102 ) ;
assign n104 =  ( n37 ) ? ( LB2D_shift_2 ) : ( LB2D_shift_2 ) ;
assign n105 =  ( n32 ) ? ( LB2D_shift_2 ) : ( n104 ) ;
assign n106 =  ( n25 ) ? ( LB2D_shift_1 ) : ( n105 ) ;
assign n107 =  ( n18 ) ? ( LB2D_shift_2 ) : ( n106 ) ;
assign n108 =  ( n9 ) ? ( LB2D_shift_2 ) : ( n107 ) ;
assign n109 =  ( n4 ) ? ( LB2D_shift_2 ) : ( n108 ) ;
assign n110 =  ( n37 ) ? ( LB2D_shift_3 ) : ( LB2D_shift_3 ) ;
assign n111 =  ( n32 ) ? ( LB2D_shift_3 ) : ( n110 ) ;
assign n112 =  ( n25 ) ? ( LB2D_shift_2 ) : ( n111 ) ;
assign n113 =  ( n18 ) ? ( LB2D_shift_3 ) : ( n112 ) ;
assign n114 =  ( n9 ) ? ( LB2D_shift_3 ) : ( n113 ) ;
assign n115 =  ( n4 ) ? ( LB2D_shift_3 ) : ( n114 ) ;
assign n116 =  ( n37 ) ? ( LB2D_shift_4 ) : ( LB2D_shift_4 ) ;
assign n117 =  ( n32 ) ? ( LB2D_shift_4 ) : ( n116 ) ;
assign n118 =  ( n25 ) ? ( LB2D_shift_3 ) : ( n117 ) ;
assign n119 =  ( n18 ) ? ( LB2D_shift_4 ) : ( n118 ) ;
assign n120 =  ( n9 ) ? ( LB2D_shift_4 ) : ( n119 ) ;
assign n121 =  ( n4 ) ? ( LB2D_shift_4 ) : ( n120 ) ;
assign n122 =  ( n37 ) ? ( LB2D_shift_5 ) : ( LB2D_shift_5 ) ;
assign n123 =  ( n32 ) ? ( LB2D_shift_5 ) : ( n122 ) ;
assign n124 =  ( n25 ) ? ( LB2D_shift_4 ) : ( n123 ) ;
assign n125 =  ( n18 ) ? ( LB2D_shift_5 ) : ( n124 ) ;
assign n126 =  ( n9 ) ? ( LB2D_shift_5 ) : ( n125 ) ;
assign n127 =  ( n4 ) ? ( LB2D_shift_5 ) : ( n126 ) ;
assign n128 =  ( n37 ) ? ( LB2D_shift_6 ) : ( LB2D_shift_6 ) ;
assign n129 =  ( n32 ) ? ( LB2D_shift_6 ) : ( n128 ) ;
assign n130 =  ( n25 ) ? ( LB2D_shift_5 ) : ( n129 ) ;
assign n131 =  ( n18 ) ? ( LB2D_shift_6 ) : ( n130 ) ;
assign n132 =  ( n9 ) ? ( LB2D_shift_6 ) : ( n131 ) ;
assign n133 =  ( n4 ) ? ( LB2D_shift_6 ) : ( n132 ) ;
assign n134 =  ( n37 ) ? ( LB2D_shift_7 ) : ( LB2D_shift_7 ) ;
assign n135 =  ( n32 ) ? ( LB2D_shift_7 ) : ( n134 ) ;
assign n136 =  ( n25 ) ? ( LB2D_shift_6 ) : ( n135 ) ;
assign n137 =  ( n18 ) ? ( LB2D_shift_7 ) : ( n136 ) ;
assign n138 =  ( n9 ) ? ( LB2D_shift_7 ) : ( n137 ) ;
assign n139 =  ( n4 ) ? ( LB2D_shift_7 ) : ( n138 ) ;
assign n140 =  ( LB2D_shift_x ) + ( 9'd1 )  ;
assign n141 =  ( n37 ) ? ( LB2D_shift_x ) : ( LB2D_shift_x ) ;
assign n142 =  ( n32 ) ? ( LB2D_shift_x ) : ( n141 ) ;
assign n143 =  ( n25 ) ? ( n140 ) : ( n142 ) ;
assign n144 =  ( n18 ) ? ( LB2D_shift_x ) : ( n143 ) ;
assign n145 =  ( n9 ) ? ( LB2D_shift_x ) : ( n144 ) ;
assign n146 =  ( n4 ) ? ( LB2D_shift_x ) : ( n145 ) ;
assign n147 =  ( LB2D_shift_y ) < ( 10'd480 )  ;
assign n148 =  ( LB2D_shift_x ) < ( 9'd488 )  ;
assign n149 =  ( LB2D_shift_y ) + ( 10'd1 )  ;
assign n150 =  ( n148 ) ? ( LB2D_shift_y ) : ( n149 ) ;
assign n151 =  ( n147 ) ? ( n150 ) : ( 10'd480 ) ;
assign n152 =  ( n37 ) ? ( LB2D_shift_y ) : ( LB2D_shift_y ) ;
assign n153 =  ( n32 ) ? ( LB2D_shift_y ) : ( n152 ) ;
assign n154 =  ( n25 ) ? ( n151 ) : ( n153 ) ;
assign n155 =  ( n18 ) ? ( LB2D_shift_y ) : ( n154 ) ;
assign n156 =  ( n9 ) ? ( LB2D_shift_y ) : ( n155 ) ;
assign n157 =  ( n4 ) ? ( LB2D_shift_y ) : ( n156 ) ;
assign n158 =  ( stencil_stream_full ) == ( 1'd1 )  ;
assign n159 =  ( n158 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_0 ) ;
//assign n160 = gb_fun(n159) ;
gb_fun gb_fun_U (
        .stencil (n159),
        .result (n160)
        );

assign n161 =  ( n37 ) ? ( arg_0_TDATA ) : ( arg_0_TDATA ) ;
assign n162 =  ( n32 ) ? ( arg_0_TDATA ) : ( n161 ) ;
assign n163 =  ( n25 ) ? ( arg_0_TDATA ) : ( n162 ) ;
assign n164 =  ( n18 ) ? ( n160 ) : ( n163 ) ;
assign n165 =  ( n9 ) ? ( arg_0_TDATA ) : ( n164 ) ;
assign n166 =  ( n4 ) ? ( arg_0_TDATA ) : ( n165 ) ;
assign n167 =  ( gb_pp_it_8 ) == ( 1'd1 )  ;
assign n168 =  ( n167 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n169 =  ( n37 ) ? ( arg_0_TVALID ) : ( arg_0_TVALID ) ;
assign n170 =  ( n32 ) ? ( arg_0_TVALID ) : ( n169 ) ;
assign n171 =  ( n25 ) ? ( arg_0_TVALID ) : ( n170 ) ;
assign n172 =  ( n18 ) ? ( n168 ) : ( n171 ) ;
assign n173 =  ( n9 ) ? ( arg_0_TVALID ) : ( n172 ) ;
assign n174 =  ( n4 ) ? ( 1'd0 ) : ( n173 ) ;
assign n175 =  ( n37 ) ? ( 1'd1 ) : ( arg_1_TREADY ) ;
assign n176 =  ( n47 ) ? ( 1'd1 ) : ( n175 ) ;
assign n177 =  ( n32 ) ? ( arg_1_TREADY ) : ( n176 ) ;
assign n178 =  ( n25 ) ? ( arg_1_TREADY ) : ( n177 ) ;
assign n179 =  ( n18 ) ? ( arg_1_TREADY ) : ( n178 ) ;
assign n180 =  ( n9 ) ? ( 1'd0 ) : ( n179 ) ;
assign n181 =  ( n4 ) ? ( 1'd0 ) : ( n180 ) ;
assign n182 =  ( gb_p_cnt ) + ( 19'd1 )  ;
assign n183 =  ( n182 ) == ( 19'd307200 )  ;
assign n184 =  ( n183 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n185 =  ( n37 ) ? ( gb_exit_it_1 ) : ( gb_exit_it_1 ) ;
assign n186 =  ( n32 ) ? ( gb_exit_it_1 ) : ( n185 ) ;
assign n187 =  ( n25 ) ? ( gb_exit_it_1 ) : ( n186 ) ;
assign n188 =  ( n18 ) ? ( n184 ) : ( n187 ) ;
assign n189 =  ( n9 ) ? ( gb_exit_it_1 ) : ( n188 ) ;
assign n190 =  ( n4 ) ? ( gb_exit_it_1 ) : ( n189 ) ;
assign n191 =  ( n37 ) ? ( gb_exit_it_2 ) : ( gb_exit_it_2 ) ;
assign n192 =  ( n32 ) ? ( gb_exit_it_2 ) : ( n191 ) ;
assign n193 =  ( n25 ) ? ( gb_exit_it_2 ) : ( n192 ) ;
assign n194 =  ( n18 ) ? ( gb_exit_it_1 ) : ( n193 ) ;
assign n195 =  ( n9 ) ? ( gb_exit_it_2 ) : ( n194 ) ;
assign n196 =  ( n4 ) ? ( gb_exit_it_2 ) : ( n195 ) ;
assign n197 =  ( n37 ) ? ( gb_exit_it_3 ) : ( gb_exit_it_3 ) ;
assign n198 =  ( n32 ) ? ( gb_exit_it_3 ) : ( n197 ) ;
assign n199 =  ( n25 ) ? ( gb_exit_it_3 ) : ( n198 ) ;
assign n200 =  ( n18 ) ? ( gb_exit_it_2 ) : ( n199 ) ;
assign n201 =  ( n9 ) ? ( gb_exit_it_3 ) : ( n200 ) ;
assign n202 =  ( n4 ) ? ( gb_exit_it_3 ) : ( n201 ) ;
assign n203 =  ( n37 ) ? ( gb_exit_it_4 ) : ( gb_exit_it_4 ) ;
assign n204 =  ( n32 ) ? ( gb_exit_it_4 ) : ( n203 ) ;
assign n205 =  ( n25 ) ? ( gb_exit_it_4 ) : ( n204 ) ;
assign n206 =  ( n18 ) ? ( gb_exit_it_3 ) : ( n205 ) ;
assign n207 =  ( n9 ) ? ( gb_exit_it_4 ) : ( n206 ) ;
assign n208 =  ( n4 ) ? ( gb_exit_it_4 ) : ( n207 ) ;
assign n209 =  ( n37 ) ? ( gb_exit_it_5 ) : ( gb_exit_it_5 ) ;
assign n210 =  ( n32 ) ? ( gb_exit_it_5 ) : ( n209 ) ;
assign n211 =  ( n25 ) ? ( gb_exit_it_5 ) : ( n210 ) ;
assign n212 =  ( n18 ) ? ( gb_exit_it_4 ) : ( n211 ) ;
assign n213 =  ( n9 ) ? ( gb_exit_it_5 ) : ( n212 ) ;
assign n214 =  ( n4 ) ? ( gb_exit_it_5 ) : ( n213 ) ;
assign n215 =  ( n37 ) ? ( gb_exit_it_6 ) : ( gb_exit_it_6 ) ;
assign n216 =  ( n32 ) ? ( gb_exit_it_6 ) : ( n215 ) ;
assign n217 =  ( n25 ) ? ( gb_exit_it_6 ) : ( n216 ) ;
assign n218 =  ( n18 ) ? ( gb_exit_it_5 ) : ( n217 ) ;
assign n219 =  ( n9 ) ? ( gb_exit_it_6 ) : ( n218 ) ;
assign n220 =  ( n4 ) ? ( gb_exit_it_6 ) : ( n219 ) ;
assign n221 =  ( n37 ) ? ( gb_exit_it_7 ) : ( gb_exit_it_7 ) ;
assign n222 =  ( n32 ) ? ( gb_exit_it_7 ) : ( n221 ) ;
assign n223 =  ( n25 ) ? ( gb_exit_it_7 ) : ( n222 ) ;
assign n224 =  ( n18 ) ? ( gb_exit_it_6 ) : ( n223 ) ;
assign n225 =  ( n9 ) ? ( gb_exit_it_7 ) : ( n224 ) ;
assign n226 =  ( n4 ) ? ( gb_exit_it_7 ) : ( n225 ) ;
assign n227 =  ( n37 ) ? ( gb_exit_it_8 ) : ( gb_exit_it_8 ) ;
assign n228 =  ( n32 ) ? ( gb_exit_it_8 ) : ( n227 ) ;
assign n229 =  ( n25 ) ? ( gb_exit_it_8 ) : ( n228 ) ;
assign n230 =  ( n18 ) ? ( gb_exit_it_7 ) : ( n229 ) ;
assign n231 =  ( n9 ) ? ( gb_exit_it_8 ) : ( n230 ) ;
assign n232 =  ( n4 ) ? ( gb_exit_it_8 ) : ( n231 ) ;
assign n233 =  ( gb_p_cnt ) < ( 19'd307200 )  ;
assign n234 =  ( n233 ) ? ( n182 ) : ( 19'd307200 ) ;
assign n235 =  ( n37 ) ? ( gb_p_cnt ) : ( gb_p_cnt ) ;
assign n236 =  ( n32 ) ? ( gb_p_cnt ) : ( n235 ) ;
assign n237 =  ( n25 ) ? ( gb_p_cnt ) : ( n236 ) ;
assign n238 =  ( n18 ) ? ( n234 ) : ( n237 ) ;
assign n239 =  ( n9 ) ? ( gb_p_cnt ) : ( n238 ) ;
assign n240 =  ( n4 ) ? ( gb_p_cnt ) : ( n239 ) ;
assign n241 =  ( n37 ) ? ( gb_pp_it_1 ) : ( gb_pp_it_1 ) ;
assign n242 =  ( n32 ) ? ( gb_pp_it_1 ) : ( n241 ) ;
assign n243 =  ( n25 ) ? ( gb_pp_it_1 ) : ( n242 ) ;
assign n244 =  ( n18 ) ? ( 1'd1 ) : ( n243 ) ;
assign n245 =  ( n9 ) ? ( gb_pp_it_1 ) : ( n244 ) ;
assign n246 =  ( n4 ) ? ( gb_pp_it_1 ) : ( n245 ) ;
assign n247 =  ( n37 ) ? ( gb_pp_it_2 ) : ( gb_pp_it_2 ) ;
assign n248 =  ( n32 ) ? ( gb_pp_it_2 ) : ( n247 ) ;
assign n249 =  ( n25 ) ? ( gb_pp_it_2 ) : ( n248 ) ;
assign n250 =  ( n18 ) ? ( gb_pp_it_1 ) : ( n249 ) ;
assign n251 =  ( n9 ) ? ( gb_pp_it_2 ) : ( n250 ) ;
assign n252 =  ( n4 ) ? ( gb_pp_it_2 ) : ( n251 ) ;
assign n253 =  ( n37 ) ? ( gb_pp_it_3 ) : ( gb_pp_it_3 ) ;
assign n254 =  ( n32 ) ? ( gb_pp_it_3 ) : ( n253 ) ;
assign n255 =  ( n25 ) ? ( gb_pp_it_3 ) : ( n254 ) ;
assign n256 =  ( n18 ) ? ( gb_pp_it_2 ) : ( n255 ) ;
assign n257 =  ( n9 ) ? ( gb_pp_it_3 ) : ( n256 ) ;
assign n258 =  ( n4 ) ? ( gb_pp_it_3 ) : ( n257 ) ;
assign n259 =  ( n37 ) ? ( gb_pp_it_4 ) : ( gb_pp_it_4 ) ;
assign n260 =  ( n32 ) ? ( gb_pp_it_4 ) : ( n259 ) ;
assign n261 =  ( n25 ) ? ( gb_pp_it_4 ) : ( n260 ) ;
assign n262 =  ( n18 ) ? ( gb_pp_it_3 ) : ( n261 ) ;
assign n263 =  ( n9 ) ? ( gb_pp_it_4 ) : ( n262 ) ;
assign n264 =  ( n4 ) ? ( gb_pp_it_4 ) : ( n263 ) ;
assign n265 =  ( n37 ) ? ( gb_pp_it_5 ) : ( gb_pp_it_5 ) ;
assign n266 =  ( n32 ) ? ( gb_pp_it_5 ) : ( n265 ) ;
assign n267 =  ( n25 ) ? ( gb_pp_it_5 ) : ( n266 ) ;
assign n268 =  ( n18 ) ? ( gb_pp_it_4 ) : ( n267 ) ;
assign n269 =  ( n9 ) ? ( gb_pp_it_5 ) : ( n268 ) ;
assign n270 =  ( n4 ) ? ( gb_pp_it_5 ) : ( n269 ) ;
assign n271 =  ( n37 ) ? ( gb_pp_it_6 ) : ( gb_pp_it_6 ) ;
assign n272 =  ( n32 ) ? ( gb_pp_it_6 ) : ( n271 ) ;
assign n273 =  ( n25 ) ? ( gb_pp_it_6 ) : ( n272 ) ;
assign n274 =  ( n18 ) ? ( gb_pp_it_5 ) : ( n273 ) ;
assign n275 =  ( n9 ) ? ( gb_pp_it_6 ) : ( n274 ) ;
assign n276 =  ( n4 ) ? ( gb_pp_it_6 ) : ( n275 ) ;
assign n277 =  ( n37 ) ? ( gb_pp_it_7 ) : ( gb_pp_it_7 ) ;
assign n278 =  ( n32 ) ? ( gb_pp_it_7 ) : ( n277 ) ;
assign n279 =  ( n25 ) ? ( gb_pp_it_7 ) : ( n278 ) ;
assign n280 =  ( n18 ) ? ( gb_pp_it_6 ) : ( n279 ) ;
assign n281 =  ( n9 ) ? ( gb_pp_it_7 ) : ( n280 ) ;
assign n282 =  ( n4 ) ? ( gb_pp_it_7 ) : ( n281 ) ;
assign n283 =  ( n37 ) ? ( gb_pp_it_8 ) : ( gb_pp_it_8 ) ;
assign n284 =  ( n32 ) ? ( gb_pp_it_8 ) : ( n283 ) ;
assign n285 =  ( n25 ) ? ( gb_pp_it_8 ) : ( n284 ) ;
assign n286 =  ( n18 ) ? ( gb_pp_it_7 ) : ( n285 ) ;
assign n287 =  ( n9 ) ? ( gb_pp_it_8 ) : ( n286 ) ;
assign n288 =  ( n4 ) ? ( gb_pp_it_8 ) : ( n287 ) ;
assign n289 =  ( n37 ) ? ( gb_pp_it_9 ) : ( gb_pp_it_9 ) ;
assign n290 =  ( n32 ) ? ( gb_pp_it_9 ) : ( n289 ) ;
assign n291 =  ( n25 ) ? ( gb_pp_it_9 ) : ( n290 ) ;
assign n292 =  ( n18 ) ? ( gb_pp_it_8 ) : ( n291 ) ;
assign n293 =  ( n9 ) ? ( gb_pp_it_9 ) : ( n292 ) ;
assign n294 =  ( n4 ) ? ( gb_pp_it_9 ) : ( n293 ) ;
assign n295 =  ( n37 ) ? ( LB1D_buff ) : ( in_stream_buff_0 ) ;
assign n296 =  ( n32 ) ? ( in_stream_buff_0 ) : ( n295 ) ;
assign n297 =  ( n25 ) ? ( in_stream_buff_0 ) : ( n296 ) ;
assign n298 =  ( n18 ) ? ( in_stream_buff_0 ) : ( n297 ) ;
assign n299 =  ( n9 ) ? ( in_stream_buff_0 ) : ( n298 ) ;
assign n300 =  ( n4 ) ? ( in_stream_buff_0 ) : ( n299 ) ;
assign n301 =  ( n37 ) ? ( in_stream_buff_0 ) : ( in_stream_buff_1 ) ;
assign n302 =  ( n32 ) ? ( in_stream_buff_1 ) : ( n301 ) ;
assign n303 =  ( n25 ) ? ( in_stream_buff_1 ) : ( n302 ) ;
assign n304 =  ( n18 ) ? ( in_stream_buff_1 ) : ( n303 ) ;
assign n305 =  ( n9 ) ? ( in_stream_buff_1 ) : ( n304 ) ;
assign n306 =  ( n4 ) ? ( in_stream_buff_1 ) : ( n305 ) ;
assign n307 =  ( in_stream_full ) == ( 1'd1 )  ;
assign n308 =  ( n307 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n309 =  ( n37 ) ? ( 1'd0 ) : ( in_stream_empty ) ;
assign n310 =  ( n32 ) ? ( n308 ) : ( n309 ) ;
assign n311 =  ( n25 ) ? ( in_stream_empty ) : ( n310 ) ;
assign n312 =  ( n18 ) ? ( in_stream_empty ) : ( n311 ) ;
assign n313 =  ( n9 ) ? ( in_stream_empty ) : ( n312 ) ;
assign n314 =  ( n4 ) ? ( in_stream_empty ) : ( n313 ) ;
assign n315 =  ( in_stream_empty ) == ( 1'd1 )  ;
assign n316 =  ( n315 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n317 =  ( n37 ) ? ( n316 ) : ( in_stream_full ) ;
assign n318 =  ( n32 ) ? ( 1'd0 ) : ( n317 ) ;
assign n319 =  ( n25 ) ? ( in_stream_full ) : ( n318 ) ;
assign n320 =  ( n18 ) ? ( in_stream_full ) : ( n319 ) ;
assign n321 =  ( n9 ) ? ( in_stream_full ) : ( n320 ) ;
assign n322 =  ( n4 ) ? ( in_stream_full ) : ( n321 ) ;
assign n323 =  ( n307 ) ? ( in_stream_buff_1 ) : ( in_stream_buff_0 ) ;
assign n324 =  ( LB2D_proc_w ) == ( 64'd0 )  ;
assign n325 =  (  LB2D_proc_7 [ LB2D_proc_x ] )  ;
assign n326 =  ( LB2D_proc_w ) == ( 64'd1 )  ;
assign n327 =  (  LB2D_proc_0 [ LB2D_proc_x ] )  ;
assign n328 =  ( LB2D_proc_w ) == ( 64'd2 )  ;
assign n329 =  (  LB2D_proc_1 [ LB2D_proc_x ] )  ;
assign n330 =  ( LB2D_proc_w ) == ( 64'd3 )  ;
assign n331 =  (  LB2D_proc_2 [ LB2D_proc_x ] )  ;
assign n332 =  ( LB2D_proc_w ) == ( 64'd4 )  ;
assign n333 =  (  LB2D_proc_3 [ LB2D_proc_x ] )  ;
assign n334 =  ( LB2D_proc_w ) == ( 64'd5 )  ;
assign n335 =  (  LB2D_proc_4 [ LB2D_proc_x ] )  ;
assign n336 =  ( LB2D_proc_w ) == ( 64'd6 )  ;
assign n337 =  (  LB2D_proc_5 [ LB2D_proc_x ] )  ;
assign n338 =  (  LB2D_proc_6 [ LB2D_proc_x ] )  ;
assign n339 =  ( n336 ) ? ( n337 ) : ( n338 ) ;
assign n340 =  ( n334 ) ? ( n335 ) : ( n339 ) ;
assign n341 =  ( n332 ) ? ( n333 ) : ( n340 ) ;
assign n342 =  ( n330 ) ? ( n331 ) : ( n341 ) ;
assign n343 =  ( n328 ) ? ( n329 ) : ( n342 ) ;
assign n344 =  ( n326 ) ? ( n327 ) : ( n343 ) ;
assign n345 =  ( n324 ) ? ( n325 ) : ( n344 ) ;
assign n346 =  ( n336 ) ? ( n335 ) : ( n337 ) ;
assign n347 =  ( n334 ) ? ( n333 ) : ( n346 ) ;
assign n348 =  ( n332 ) ? ( n331 ) : ( n347 ) ;
assign n349 =  ( n330 ) ? ( n329 ) : ( n348 ) ;
assign n350 =  ( n328 ) ? ( n327 ) : ( n349 ) ;
assign n351 =  ( n326 ) ? ( n325 ) : ( n350 ) ;
assign n352 =  ( n324 ) ? ( n338 ) : ( n351 ) ;
assign n353 =  ( n336 ) ? ( n333 ) : ( n335 ) ;
assign n354 =  ( n334 ) ? ( n331 ) : ( n353 ) ;
assign n355 =  ( n332 ) ? ( n329 ) : ( n354 ) ;
assign n356 =  ( n330 ) ? ( n327 ) : ( n355 ) ;
assign n357 =  ( n328 ) ? ( n325 ) : ( n356 ) ;
assign n358 =  ( n326 ) ? ( n338 ) : ( n357 ) ;
assign n359 =  ( n324 ) ? ( n337 ) : ( n358 ) ;
assign n360 =  ( n336 ) ? ( n331 ) : ( n333 ) ;
assign n361 =  ( n334 ) ? ( n329 ) : ( n360 ) ;
assign n362 =  ( n332 ) ? ( n327 ) : ( n361 ) ;
assign n363 =  ( n330 ) ? ( n325 ) : ( n362 ) ;
assign n364 =  ( n328 ) ? ( n338 ) : ( n363 ) ;
assign n365 =  ( n326 ) ? ( n337 ) : ( n364 ) ;
assign n366 =  ( n324 ) ? ( n335 ) : ( n365 ) ;
assign n367 =  ( n336 ) ? ( n329 ) : ( n331 ) ;
assign n368 =  ( n334 ) ? ( n327 ) : ( n367 ) ;
assign n369 =  ( n332 ) ? ( n325 ) : ( n368 ) ;
assign n370 =  ( n330 ) ? ( n338 ) : ( n369 ) ;
assign n371 =  ( n328 ) ? ( n337 ) : ( n370 ) ;
assign n372 =  ( n326 ) ? ( n335 ) : ( n371 ) ;
assign n373 =  ( n324 ) ? ( n333 ) : ( n372 ) ;
assign n374 =  ( n336 ) ? ( n327 ) : ( n329 ) ;
assign n375 =  ( n334 ) ? ( n325 ) : ( n374 ) ;
assign n376 =  ( n332 ) ? ( n338 ) : ( n375 ) ;
assign n377 =  ( n330 ) ? ( n337 ) : ( n376 ) ;
assign n378 =  ( n328 ) ? ( n335 ) : ( n377 ) ;
assign n379 =  ( n326 ) ? ( n333 ) : ( n378 ) ;
assign n380 =  ( n324 ) ? ( n331 ) : ( n379 ) ;
assign n381 =  ( n336 ) ? ( n325 ) : ( n327 ) ;
assign n382 =  ( n334 ) ? ( n338 ) : ( n381 ) ;
assign n383 =  ( n332 ) ? ( n337 ) : ( n382 ) ;
assign n384 =  ( n330 ) ? ( n335 ) : ( n383 ) ;
assign n385 =  ( n328 ) ? ( n333 ) : ( n384 ) ;
assign n386 =  ( n326 ) ? ( n331 ) : ( n385 ) ;
assign n387 =  ( n324 ) ? ( n329 ) : ( n386 ) ;
assign n388 =  ( n336 ) ? ( n338 ) : ( n325 ) ;
assign n389 =  ( n334 ) ? ( n337 ) : ( n388 ) ;
assign n390 =  ( n332 ) ? ( n335 ) : ( n389 ) ;
assign n391 =  ( n330 ) ? ( n333 ) : ( n390 ) ;
assign n392 =  ( n328 ) ? ( n331 ) : ( n391 ) ;
assign n393 =  ( n326 ) ? ( n329 ) : ( n392 ) ;
assign n394 =  ( n324 ) ? ( n327 ) : ( n393 ) ;
assign n395 =  { ( n387 ) , ( n394 ) }  ;
assign n396 =  { ( n380 ) , ( n395 ) }  ;
assign n397 =  { ( n373 ) , ( n396 ) }  ;
assign n398 =  { ( n366 ) , ( n397 ) }  ;
assign n399 =  { ( n359 ) , ( n398 ) }  ;
assign n400 =  { ( n352 ) , ( n399 ) }  ;
assign n401 =  { ( n345 ) , ( n400 ) }  ;
assign n402 =  { ( n323 ) , ( n401 ) }  ;
assign n403 =  ( n30 ) ? ( slice_stream_buff_0 ) : ( n402 ) ;
assign n404 =  ( n37 ) ? ( slice_stream_buff_0 ) : ( slice_stream_buff_0 ) ;
assign n405 =  ( n32 ) ? ( n403 ) : ( n404 ) ;
assign n406 =  ( n25 ) ? ( slice_stream_buff_0 ) : ( n405 ) ;
assign n407 =  ( n18 ) ? ( slice_stream_buff_0 ) : ( n406 ) ;
assign n408 =  ( n9 ) ? ( slice_stream_buff_0 ) : ( n407 ) ;
assign n409 =  ( n4 ) ? ( slice_stream_buff_0 ) : ( n408 ) ;
assign n410 =  ( n30 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n411 =  ( n37 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_1 ) ;
assign n412 =  ( n32 ) ? ( n410 ) : ( n411 ) ;
assign n413 =  ( n25 ) ? ( slice_stream_buff_1 ) : ( n412 ) ;
assign n414 =  ( n18 ) ? ( slice_stream_buff_1 ) : ( n413 ) ;
assign n415 =  ( n9 ) ? ( slice_stream_buff_1 ) : ( n414 ) ;
assign n416 =  ( n4 ) ? ( slice_stream_buff_1 ) : ( n415 ) ;
assign n417 =  ( n90 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n418 =  ( n30 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n419 =  ( n37 ) ? ( slice_stream_empty ) : ( slice_stream_empty ) ;
assign n420 =  ( n32 ) ? ( n418 ) : ( n419 ) ;
assign n421 =  ( n25 ) ? ( n417 ) : ( n420 ) ;
assign n422 =  ( n18 ) ? ( slice_stream_empty ) : ( n421 ) ;
assign n423 =  ( n9 ) ? ( slice_stream_empty ) : ( n422 ) ;
assign n424 =  ( n4 ) ? ( slice_stream_empty ) : ( n423 ) ;
assign n425 =  ( slice_stream_empty ) == ( 1'd1 )  ;
assign n426 =  ( n425 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n427 =  ( n30 ) ? ( 1'd0 ) : ( n426 ) ;
assign n428 =  ( n37 ) ? ( slice_stream_full ) : ( slice_stream_full ) ;
assign n429 =  ( n32 ) ? ( n427 ) : ( n428 ) ;
assign n430 =  ( n25 ) ? ( 1'd0 ) : ( n429 ) ;
assign n431 =  ( n18 ) ? ( slice_stream_full ) : ( n430 ) ;
assign n432 =  ( n9 ) ? ( slice_stream_full ) : ( n431 ) ;
assign n433 =  ( n4 ) ? ( slice_stream_full ) : ( n432 ) ;
assign n434 =  ( LB2D_shift_x ) >= ( 9'd8 )  ;
assign n435 = n91[71:64] ;
assign n436 = LB2D_shift_0[71:64] ;
assign n437 = LB2D_shift_1[71:64] ;
assign n438 = LB2D_shift_2[71:64] ;
assign n439 = LB2D_shift_3[71:64] ;
assign n440 = LB2D_shift_4[71:64] ;
assign n441 = LB2D_shift_5[71:64] ;
assign n442 = LB2D_shift_6[71:64] ;
assign n443 = LB2D_shift_7[71:64] ;
assign n444 =  { ( n442 ) , ( n443 ) }  ;
assign n445 =  { ( n441 ) , ( n444 ) }  ;
assign n446 =  { ( n440 ) , ( n445 ) }  ;
assign n447 =  { ( n439 ) , ( n446 ) }  ;
assign n448 =  { ( n438 ) , ( n447 ) }  ;
assign n449 =  { ( n437 ) , ( n448 ) }  ;
assign n450 =  { ( n436 ) , ( n449 ) }  ;
assign n451 =  { ( n435 ) , ( n450 ) }  ;
assign n452 = n91[63:56] ;
assign n453 = LB2D_shift_0[63:56] ;
assign n454 = LB2D_shift_1[63:56] ;
assign n455 = LB2D_shift_2[63:56] ;
assign n456 = LB2D_shift_3[63:56] ;
assign n457 = LB2D_shift_4[63:56] ;
assign n458 = LB2D_shift_5[63:56] ;
assign n459 = LB2D_shift_6[63:56] ;
assign n460 = LB2D_shift_7[63:56] ;
assign n461 =  { ( n459 ) , ( n460 ) }  ;
assign n462 =  { ( n458 ) , ( n461 ) }  ;
assign n463 =  { ( n457 ) , ( n462 ) }  ;
assign n464 =  { ( n456 ) , ( n463 ) }  ;
assign n465 =  { ( n455 ) , ( n464 ) }  ;
assign n466 =  { ( n454 ) , ( n465 ) }  ;
assign n467 =  { ( n453 ) , ( n466 ) }  ;
assign n468 =  { ( n452 ) , ( n467 ) }  ;
assign n469 = n91[55:48] ;
assign n470 = LB2D_shift_0[55:48] ;
assign n471 = LB2D_shift_1[55:48] ;
assign n472 = LB2D_shift_2[55:48] ;
assign n473 = LB2D_shift_3[55:48] ;
assign n474 = LB2D_shift_4[55:48] ;
assign n475 = LB2D_shift_5[55:48] ;
assign n476 = LB2D_shift_6[55:48] ;
assign n477 = LB2D_shift_7[55:48] ;
assign n478 =  { ( n476 ) , ( n477 ) }  ;
assign n479 =  { ( n475 ) , ( n478 ) }  ;
assign n480 =  { ( n474 ) , ( n479 ) }  ;
assign n481 =  { ( n473 ) , ( n480 ) }  ;
assign n482 =  { ( n472 ) , ( n481 ) }  ;
assign n483 =  { ( n471 ) , ( n482 ) }  ;
assign n484 =  { ( n470 ) , ( n483 ) }  ;
assign n485 =  { ( n469 ) , ( n484 ) }  ;
assign n486 = n91[47:40] ;
assign n487 = LB2D_shift_0[47:40] ;
assign n488 = LB2D_shift_1[47:40] ;
assign n489 = LB2D_shift_2[47:40] ;
assign n490 = LB2D_shift_3[47:40] ;
assign n491 = LB2D_shift_4[47:40] ;
assign n492 = LB2D_shift_5[47:40] ;
assign n493 = LB2D_shift_6[47:40] ;
assign n494 = LB2D_shift_7[47:40] ;
assign n495 =  { ( n493 ) , ( n494 ) }  ;
assign n496 =  { ( n492 ) , ( n495 ) }  ;
assign n497 =  { ( n491 ) , ( n496 ) }  ;
assign n498 =  { ( n490 ) , ( n497 ) }  ;
assign n499 =  { ( n489 ) , ( n498 ) }  ;
assign n500 =  { ( n488 ) , ( n499 ) }  ;
assign n501 =  { ( n487 ) , ( n500 ) }  ;
assign n502 =  { ( n486 ) , ( n501 ) }  ;
assign n503 = n91[39:32] ;
assign n504 = LB2D_shift_0[39:32] ;
assign n505 = LB2D_shift_1[39:32] ;
assign n506 = LB2D_shift_2[39:32] ;
assign n507 = LB2D_shift_3[39:32] ;
assign n508 = LB2D_shift_4[39:32] ;
assign n509 = LB2D_shift_5[39:32] ;
assign n510 = LB2D_shift_6[39:32] ;
assign n511 = LB2D_shift_7[39:32] ;
assign n512 =  { ( n510 ) , ( n511 ) }  ;
assign n513 =  { ( n509 ) , ( n512 ) }  ;
assign n514 =  { ( n508 ) , ( n513 ) }  ;
assign n515 =  { ( n507 ) , ( n514 ) }  ;
assign n516 =  { ( n506 ) , ( n515 ) }  ;
assign n517 =  { ( n505 ) , ( n516 ) }  ;
assign n518 =  { ( n504 ) , ( n517 ) }  ;
assign n519 =  { ( n503 ) , ( n518 ) }  ;
assign n520 = n91[31:24] ;
assign n521 = LB2D_shift_0[31:24] ;
assign n522 = LB2D_shift_1[31:24] ;
assign n523 = LB2D_shift_2[31:24] ;
assign n524 = LB2D_shift_3[31:24] ;
assign n525 = LB2D_shift_4[31:24] ;
assign n526 = LB2D_shift_5[31:24] ;
assign n527 = LB2D_shift_6[31:24] ;
assign n528 = LB2D_shift_7[31:24] ;
assign n529 =  { ( n527 ) , ( n528 ) }  ;
assign n530 =  { ( n526 ) , ( n529 ) }  ;
assign n531 =  { ( n525 ) , ( n530 ) }  ;
assign n532 =  { ( n524 ) , ( n531 ) }  ;
assign n533 =  { ( n523 ) , ( n532 ) }  ;
assign n534 =  { ( n522 ) , ( n533 ) }  ;
assign n535 =  { ( n521 ) , ( n534 ) }  ;
assign n536 =  { ( n520 ) , ( n535 ) }  ;
assign n537 = n91[23:16] ;
assign n538 = LB2D_shift_0[23:16] ;
assign n539 = LB2D_shift_1[23:16] ;
assign n540 = LB2D_shift_2[23:16] ;
assign n541 = LB2D_shift_3[23:16] ;
assign n542 = LB2D_shift_4[23:16] ;
assign n543 = LB2D_shift_5[23:16] ;
assign n544 = LB2D_shift_6[23:16] ;
assign n545 = LB2D_shift_7[23:16] ;
assign n546 =  { ( n544 ) , ( n545 ) }  ;
assign n547 =  { ( n543 ) , ( n546 ) }  ;
assign n548 =  { ( n542 ) , ( n547 ) }  ;
assign n549 =  { ( n541 ) , ( n548 ) }  ;
assign n550 =  { ( n540 ) , ( n549 ) }  ;
assign n551 =  { ( n539 ) , ( n550 ) }  ;
assign n552 =  { ( n538 ) , ( n551 ) }  ;
assign n553 =  { ( n537 ) , ( n552 ) }  ;
assign n554 = n91[15:8] ;
assign n555 = LB2D_shift_0[15:8] ;
assign n556 = LB2D_shift_1[15:8] ;
assign n557 = LB2D_shift_2[15:8] ;
assign n558 = LB2D_shift_3[15:8] ;
assign n559 = LB2D_shift_4[15:8] ;
assign n560 = LB2D_shift_5[15:8] ;
assign n561 = LB2D_shift_6[15:8] ;
assign n562 = LB2D_shift_7[15:8] ;
assign n563 =  { ( n561 ) , ( n562 ) }  ;
assign n564 =  { ( n560 ) , ( n563 ) }  ;
assign n565 =  { ( n559 ) , ( n564 ) }  ;
assign n566 =  { ( n558 ) , ( n565 ) }  ;
assign n567 =  { ( n557 ) , ( n566 ) }  ;
assign n568 =  { ( n556 ) , ( n567 ) }  ;
assign n569 =  { ( n555 ) , ( n568 ) }  ;
assign n570 =  { ( n554 ) , ( n569 ) }  ;
assign n571 = n91[7:0] ;
assign n572 = LB2D_shift_0[7:0] ;
assign n573 = LB2D_shift_1[7:0] ;
assign n574 = LB2D_shift_2[7:0] ;
assign n575 = LB2D_shift_3[7:0] ;
assign n576 = LB2D_shift_4[7:0] ;
assign n577 = LB2D_shift_5[7:0] ;
assign n578 = LB2D_shift_6[7:0] ;
assign n579 = LB2D_shift_7[7:0] ;
assign n580 =  { ( n578 ) , ( n579 ) }  ;
assign n581 =  { ( n577 ) , ( n580 ) }  ;
assign n582 =  { ( n576 ) , ( n581 ) }  ;
assign n583 =  { ( n575 ) , ( n582 ) }  ;
assign n584 =  { ( n574 ) , ( n583 ) }  ;
assign n585 =  { ( n573 ) , ( n584 ) }  ;
assign n586 =  { ( n572 ) , ( n585 ) }  ;
assign n587 =  { ( n571 ) , ( n586 ) }  ;
assign n588 =  { ( n570 ) , ( n587 ) }  ;
assign n589 =  { ( n553 ) , ( n588 ) }  ;
assign n590 =  { ( n536 ) , ( n589 ) }  ;
assign n591 =  { ( n519 ) , ( n590 ) }  ;
assign n592 =  { ( n502 ) , ( n591 ) }  ;
assign n593 =  { ( n485 ) , ( n592 ) }  ;
assign n594 =  { ( n468 ) , ( n593 ) }  ;
assign n595 =  { ( n451 ) , ( n594 ) }  ;
assign n596 =  ( n434 ) ? ( n595 ) : ( stencil_stream_buff_0 ) ;
assign n597 =  ( n37 ) ? ( stencil_stream_buff_0 ) : ( stencil_stream_buff_0 ) ;
assign n598 =  ( n32 ) ? ( stencil_stream_buff_0 ) : ( n597 ) ;
assign n599 =  ( n25 ) ? ( n596 ) : ( n598 ) ;
assign n600 =  ( n18 ) ? ( stencil_stream_buff_0 ) : ( n599 ) ;
assign n601 =  ( n9 ) ? ( stencil_stream_buff_0 ) : ( n600 ) ;
assign n602 =  ( n4 ) ? ( stencil_stream_buff_0 ) : ( n601 ) ;
assign n603 =  ( n37 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_1 ) ;
assign n604 =  ( n32 ) ? ( stencil_stream_buff_1 ) : ( n603 ) ;
assign n605 =  ( n25 ) ? ( stencil_stream_buff_0 ) : ( n604 ) ;
assign n606 =  ( n18 ) ? ( stencil_stream_buff_1 ) : ( n605 ) ;
assign n607 =  ( n9 ) ? ( stencil_stream_buff_1 ) : ( n606 ) ;
assign n608 =  ( n4 ) ? ( stencil_stream_buff_1 ) : ( n607 ) ;
assign n609 =  ( n158 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n610 =  ( n23 ) ? ( stencil_stream_empty ) : ( 1'd0 ) ;
assign n611 =  ( n37 ) ? ( stencil_stream_empty ) : ( stencil_stream_empty ) ;
assign n612 =  ( n32 ) ? ( stencil_stream_empty ) : ( n611 ) ;
assign n613 =  ( n25 ) ? ( n610 ) : ( n612 ) ;
assign n614 =  ( n18 ) ? ( n609 ) : ( n613 ) ;
assign n615 =  ( n9 ) ? ( stencil_stream_empty ) : ( n614 ) ;
assign n616 =  ( n4 ) ? ( stencil_stream_empty ) : ( n615 ) ;
assign n617 =  ( n14 ) ? ( 1'd0 ) : ( 1'd0 ) ;
assign n618 =  ( stencil_stream_empty ) == ( 1'd1 )  ;
assign n619 =  ( n618 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n620 =  ( n23 ) ? ( stencil_stream_full ) : ( n619 ) ;
assign n621 =  ( n37 ) ? ( stencil_stream_full ) : ( stencil_stream_full ) ;
assign n622 =  ( n32 ) ? ( stencil_stream_full ) : ( n621 ) ;
assign n623 =  ( n25 ) ? ( n620 ) : ( n622 ) ;
assign n624 =  ( n18 ) ? ( n617 ) : ( n623 ) ;
assign n625 =  ( n9 ) ? ( stencil_stream_full ) : ( n624 ) ;
assign n626 =  ( n4 ) ? ( stencil_stream_full ) : ( n625 ) ;
assign n627 = ~ ( n4 ) ;
assign n628 = ~ ( n9 ) ;
assign n629 =  ( n627 ) & ( n628 )  ;
assign n630 = ~ ( n18 ) ;
assign n631 =  ( n629 ) & ( n630 )  ;
assign n632 = ~ ( n25 ) ;
assign n633 =  ( n631 ) & ( n632 )  ;
assign n634 = ~ ( n32 ) ;
assign n635 =  ( n633 ) & ( n634 )  ;
assign n636 = ~ ( n37 ) ;
assign n637 =  ( n635 ) & ( n636 )  ;
assign n638 =  ( n635 ) & ( n37 )  ;
assign n639 =  ( n633 ) & ( n32 )  ;
assign n640 = ~ ( n324 ) ;
assign n641 =  ( n639 ) & ( n640 )  ;
assign n642 =  ( n639 ) & ( n324 )  ;
assign n643 =  ( n631 ) & ( n25 )  ;
assign n644 =  ( n629 ) & ( n18 )  ;
assign n645 =  ( n627 ) & ( n9 )  ;
assign LB2D_proc_0_addr0 = n642 ? (LB2D_proc_x) : (0);
assign LB2D_proc_0_data0 = n642 ? (n323) : (LB2D_proc_0[0]);
assign n646 = ~ ( n326 ) ;
assign n647 =  ( n639 ) & ( n646 )  ;
assign n648 =  ( n639 ) & ( n326 )  ;
assign LB2D_proc_1_addr0 = n648 ? (LB2D_proc_x) : (0);
assign LB2D_proc_1_data0 = n648 ? (n323) : (LB2D_proc_1[0]);
assign n649 = ~ ( n328 ) ;
assign n650 =  ( n639 ) & ( n649 )  ;
assign n651 =  ( n639 ) & ( n328 )  ;
assign LB2D_proc_2_addr0 = n651 ? (LB2D_proc_x) : (0);
assign LB2D_proc_2_data0 = n651 ? (n323) : (LB2D_proc_2[0]);
assign n652 = ~ ( n330 ) ;
assign n653 =  ( n639 ) & ( n652 )  ;
assign n654 =  ( n639 ) & ( n330 )  ;
assign LB2D_proc_3_addr0 = n654 ? (LB2D_proc_x) : (0);
assign LB2D_proc_3_data0 = n654 ? (n323) : (LB2D_proc_3[0]);
assign n655 = ~ ( n332 ) ;
assign n656 =  ( n639 ) & ( n655 )  ;
assign n657 =  ( n639 ) & ( n332 )  ;
assign LB2D_proc_4_addr0 = n657 ? (LB2D_proc_x) : (0);
assign LB2D_proc_4_data0 = n657 ? (n323) : (LB2D_proc_4[0]);
assign n658 = ~ ( n334 ) ;
assign n659 =  ( n639 ) & ( n658 )  ;
assign n660 =  ( n639 ) & ( n334 )  ;
assign LB2D_proc_5_addr0 = n660 ? (LB2D_proc_x) : (0);
assign LB2D_proc_5_data0 = n660 ? (n323) : (LB2D_proc_5[0]);
assign n661 = ~ ( n336 ) ;
assign n662 =  ( n639 ) & ( n661 )  ;
assign n663 =  ( n639 ) & ( n336 )  ;
assign LB2D_proc_6_addr0 = n663 ? (LB2D_proc_x) : (0);
assign LB2D_proc_6_data0 = n663 ? (n323) : (LB2D_proc_6[0]);
assign n664 =  ( LB2D_proc_w ) == ( 64'd7 )  ;
assign n665 = ~ ( n664 ) ;
assign n666 =  ( n639 ) & ( n665 )  ;
assign n667 =  ( n639 ) & ( n664 )  ;
assign LB2D_proc_7_addr0 = n667 ? (LB2D_proc_x) : (0);
assign LB2D_proc_7_data0 = n667 ? (n323) : (LB2D_proc_7[0]);
/*
function [7:0] gb_fun ;
input [647:0] arg0;
    begin
//TODO: Add the specific function HERE.    end
endfunction
*/

always @(posedge clk) begin
   if(rst) begin
       LB1D_buff <= LB1D_buff;
       LB1D_in <= LB1D_in;
       LB1D_it_1 <= LB1D_it_1;
       LB1D_p_cnt <= LB1D_p_cnt;
       LB2D_proc_w <= LB2D_proc_w;
       LB2D_proc_x <= LB2D_proc_x;
       LB2D_proc_y <= LB2D_proc_y;
       LB2D_shift_0 <= LB2D_shift_0;
       LB2D_shift_1 <= LB2D_shift_1;
       LB2D_shift_2 <= LB2D_shift_2;
       LB2D_shift_3 <= LB2D_shift_3;
       LB2D_shift_4 <= LB2D_shift_4;
       LB2D_shift_5 <= LB2D_shift_5;
       LB2D_shift_6 <= LB2D_shift_6;
       LB2D_shift_7 <= LB2D_shift_7;
       LB2D_shift_x <= LB2D_shift_x;
       LB2D_shift_y <= LB2D_shift_y;
       arg_0_TDATA <= arg_0_TDATA;
       arg_0_TVALID <= arg_0_TVALID;
       arg_1_TREADY <= arg_1_TREADY;
       gb_exit_it_1 <= gb_exit_it_1;
       gb_exit_it_2 <= gb_exit_it_2;
       gb_exit_it_3 <= gb_exit_it_3;
       gb_exit_it_4 <= gb_exit_it_4;
       gb_exit_it_5 <= gb_exit_it_5;
       gb_exit_it_6 <= gb_exit_it_6;
       gb_exit_it_7 <= gb_exit_it_7;
       gb_exit_it_8 <= gb_exit_it_8;
       gb_p_cnt <= gb_p_cnt;
       gb_pp_it_1 <= gb_pp_it_1;
       gb_pp_it_2 <= gb_pp_it_2;
       gb_pp_it_3 <= gb_pp_it_3;
       gb_pp_it_4 <= gb_pp_it_4;
       gb_pp_it_5 <= gb_pp_it_5;
       gb_pp_it_6 <= gb_pp_it_6;
       gb_pp_it_7 <= gb_pp_it_7;
       gb_pp_it_8 <= gb_pp_it_8;
       gb_pp_it_9 <= gb_pp_it_9;
       in_stream_buff_0 <= in_stream_buff_0;
       in_stream_buff_1 <= in_stream_buff_1;
       in_stream_empty <= in_stream_empty;
       in_stream_full <= in_stream_full;
       slice_stream_buff_0 <= slice_stream_buff_0;
       slice_stream_buff_1 <= slice_stream_buff_1;
       slice_stream_empty <= slice_stream_empty;
       slice_stream_full <= slice_stream_full;
       stencil_stream_buff_0 <= stencil_stream_buff_0;
       stencil_stream_buff_1 <= stencil_stream_buff_1;
       stencil_stream_empty <= stencil_stream_empty;
       stencil_stream_full <= stencil_stream_full;
   end
   else if(step) begin
       LB1D_buff <= n43;
       LB1D_in <= n45;
       LB1D_it_1 <= n48;
       LB1D_p_cnt <= n59;
       LB2D_proc_w <= n70;
       LB2D_proc_x <= n81;
       LB2D_proc_y <= n89;
       LB2D_shift_0 <= n97;
       LB2D_shift_1 <= n103;
       LB2D_shift_2 <= n109;
       LB2D_shift_3 <= n115;
       LB2D_shift_4 <= n121;
       LB2D_shift_5 <= n127;
       LB2D_shift_6 <= n133;
       LB2D_shift_7 <= n139;
       LB2D_shift_x <= n146;
       LB2D_shift_y <= n157;
       arg_0_TDATA <= n166;
       arg_0_TVALID <= n174;
       arg_1_TREADY <= n181;
       gb_exit_it_1 <= n190;
       gb_exit_it_2 <= n196;
       gb_exit_it_3 <= n202;
       gb_exit_it_4 <= n208;
       gb_exit_it_5 <= n214;
       gb_exit_it_6 <= n220;
       gb_exit_it_7 <= n226;
       gb_exit_it_8 <= n232;
       gb_p_cnt <= n240;
       gb_pp_it_1 <= n246;
       gb_pp_it_2 <= n252;
       gb_pp_it_3 <= n258;
       gb_pp_it_4 <= n264;
       gb_pp_it_5 <= n270;
       gb_pp_it_6 <= n276;
       gb_pp_it_7 <= n282;
       gb_pp_it_8 <= n288;
       gb_pp_it_9 <= n294;
       in_stream_buff_0 <= n300;
       in_stream_buff_1 <= n306;
       in_stream_empty <= n314;
       in_stream_full <= n322;
       slice_stream_buff_0 <= n409;
       slice_stream_buff_1 <= n416;
       slice_stream_empty <= n424;
       slice_stream_full <= n433;
       stencil_stream_buff_0 <= n602;
       stencil_stream_buff_1 <= n608;
       stencil_stream_empty <= n616;
       stencil_stream_full <= n626;
       LB2D_proc_0 [ LB2D_proc_0_addr0 ] <= LB2D_proc_0_data0;
       LB2D_proc_1 [ LB2D_proc_1_addr0 ] <= LB2D_proc_1_data0;
       LB2D_proc_2 [ LB2D_proc_2_addr0 ] <= LB2D_proc_2_data0;
       LB2D_proc_3 [ LB2D_proc_3_addr0 ] <= LB2D_proc_3_data0;
       LB2D_proc_4 [ LB2D_proc_4_addr0 ] <= LB2D_proc_4_data0;
       LB2D_proc_5 [ LB2D_proc_5_addr0 ] <= LB2D_proc_5_data0;
       LB2D_proc_6 [ LB2D_proc_6_addr0 ] <= LB2D_proc_6_data0;
       LB2D_proc_7 [ LB2D_proc_7_addr0 ] <= LB2D_proc_7_data0;
   end
end
endmodule
