module GB(
arg_0_TREADY,
arg_1_TDATA,
arg_1_TVALID,
LB1D_buff,
LB2D_proc_w,
LB2D_proc_x,
LB2D_proc_y,
LB2D_shift_0,
LB2D_shift_1,
LB2D_shift_2,
LB2D_shift_3,
LB2D_shift_4,
LB2D_shift_5,
LB2D_shift_6,
LB2D_shift_7,
LB2D_shift_x,
LB2D_shift_y,
arg_0_TDATA,
arg_0_TVALID,
arg_1_TREADY,
in_stream_buff_0,
in_stream_buff_1,
in_stream_empty,
in_stream_full,
slice_stream_buff_0,
slice_stream_buff_1,
slice_stream_empty,
slice_stream_full,
stencil_stream_buff_0,
stencil_stream_buff_1,
stencil_stream_empty,
stencil_stream_full,
clk,rst,
step
);
input            arg_0_TREADY;
input      [7:0] arg_1_TDATA;
input            arg_1_TVALID;
input clk;
input rst;
input step;
output      [7:0] LB1D_buff;
output     [63:0] LB2D_proc_w;
output      [8:0] LB2D_proc_x;
output      [9:0] LB2D_proc_y;
output     [71:0] LB2D_shift_0;
output     [71:0] LB2D_shift_1;
output     [71:0] LB2D_shift_2;
output     [71:0] LB2D_shift_3;
output     [71:0] LB2D_shift_4;
output     [71:0] LB2D_shift_5;
output     [71:0] LB2D_shift_6;
output     [71:0] LB2D_shift_7;
output      [8:0] LB2D_shift_x;
output      [9:0] LB2D_shift_y;
output      [7:0] arg_0_TDATA;
output            arg_0_TVALID;
output            arg_1_TREADY;
output      [7:0] in_stream_buff_0;
output      [7:0] in_stream_buff_1;
output            in_stream_empty;
output            in_stream_full;
output     [71:0] slice_stream_buff_0;
output     [71:0] slice_stream_buff_1;
output            slice_stream_empty;
output            slice_stream_full;
output    [647:0] stencil_stream_buff_0;
output    [647:0] stencil_stream_buff_1;
output            stencil_stream_empty;
output            stencil_stream_full;
reg      [7:0] LB1D_buff;
reg     [63:0] LB2D_proc_w;
reg      [8:0] LB2D_proc_x;
reg      [9:0] LB2D_proc_y;
reg     [71:0] LB2D_shift_0;
reg     [71:0] LB2D_shift_1;
reg     [71:0] LB2D_shift_2;
reg     [71:0] LB2D_shift_3;
reg     [71:0] LB2D_shift_4;
reg     [71:0] LB2D_shift_5;
reg     [71:0] LB2D_shift_6;
reg     [71:0] LB2D_shift_7;
reg      [8:0] LB2D_shift_x;
reg      [9:0] LB2D_shift_y;
reg      [7:0] arg_0_TDATA;
reg            arg_0_TVALID;
reg            arg_1_TREADY;
reg      [7:0] in_stream_buff_0;
reg      [7:0] in_stream_buff_1;
reg            in_stream_empty;
reg            in_stream_full;
reg     [71:0] slice_stream_buff_0;
reg     [71:0] slice_stream_buff_1;
reg            slice_stream_empty;
reg            slice_stream_full;
reg    [647:0] stencil_stream_buff_0;
reg    [647:0] stencil_stream_buff_1;
reg            stencil_stream_empty;
reg            stencil_stream_full;
wire            arg_0_TREADY;
wire      [7:0] arg_1_TDATA;
wire            arg_1_TVALID;
wire            n0;
wire            n1;
wire            n2;
wire            n3;
wire            n4;
wire            n5;
wire            n6;
wire            n7;
wire            n8;
wire            n9;
wire            n10;
wire            n11;
wire            n12;
wire            n13;
wire            n14;
wire            n15;
wire            n16;
wire            n17;
wire            n18;
wire      [7:0] n19;
wire      [7:0] n20;
wire      [7:0] n21;
wire      [7:0] n22;
wire      [7:0] n23;
wire            n24;
wire            n25;
wire     [63:0] n26;
wire     [63:0] n27;
wire     [63:0] n28;
wire     [63:0] n29;
wire     [63:0] n30;
wire     [63:0] n31;
wire     [63:0] n32;
wire     [63:0] n33;
wire      [8:0] n34;
wire      [8:0] n35;
wire      [8:0] n36;
wire      [8:0] n37;
wire      [8:0] n38;
wire      [8:0] n39;
wire      [8:0] n40;
wire            n41;
wire      [9:0] n42;
wire      [9:0] n43;
wire      [9:0] n44;
wire      [9:0] n45;
wire      [9:0] n46;
wire      [9:0] n47;
wire      [9:0] n48;
wire      [9:0] n49;
wire            n50;
wire     [71:0] n51;
wire     [71:0] n52;
wire     [71:0] n53;
wire     [71:0] n54;
wire     [71:0] n55;
wire     [71:0] n56;
wire     [71:0] n57;
wire     [71:0] n58;
wire     [71:0] n59;
wire     [71:0] n60;
wire     [71:0] n61;
wire     [71:0] n62;
wire     [71:0] n63;
wire     [71:0] n64;
wire     [71:0] n65;
wire     [71:0] n66;
wire     [71:0] n67;
wire     [71:0] n68;
wire     [71:0] n69;
wire     [71:0] n70;
wire     [71:0] n71;
wire     [71:0] n72;
wire     [71:0] n73;
wire     [71:0] n74;
wire     [71:0] n75;
wire     [71:0] n76;
wire     [71:0] n77;
wire     [71:0] n78;
wire     [71:0] n79;
wire     [71:0] n80;
wire     [71:0] n81;
wire     [71:0] n82;
wire     [71:0] n83;
wire     [71:0] n84;
wire     [71:0] n85;
wire     [71:0] n86;
wire     [71:0] n87;
wire     [71:0] n88;
wire     [71:0] n89;
wire     [71:0] n90;
wire     [71:0] n91;
wire            n92;
wire      [8:0] n93;
wire      [8:0] n94;
wire      [8:0] n95;
wire      [8:0] n96;
wire      [8:0] n97;
wire      [8:0] n98;
wire      [8:0] n99;
wire      [9:0] n100;
wire      [9:0] n101;
wire      [9:0] n102;
wire      [9:0] n103;
wire      [9:0] n104;
wire      [7:0] n105;
wire      [7:0] n106;
wire      [7:0] n107;
wire      [7:0] n108;
wire      [7:0] n109;
wire            n110;
wire            n111;
wire            n112;
wire            n113;
wire            n114;
wire            n115;
wire            n116;
wire            n117;
wire            n118;
wire            n119;
wire      [7:0] n120;
wire      [7:0] n121;
wire      [7:0] n122;
wire      [7:0] n123;
wire      [7:0] n124;
wire      [7:0] n125;
wire      [7:0] n126;
wire      [7:0] n127;
wire      [7:0] n128;
wire      [7:0] n129;
wire            n130;
wire            n131;
wire            n132;
wire            n133;
wire            n134;
wire            n135;
wire            n136;
wire            n137;
wire            n138;
wire            n139;
wire            n140;
wire            n141;
wire            n142;
wire            n143;
wire            n144;
wire      [7:0] n145;
wire            n146;
wire      [7:0] n147;
wire            n148;
wire      [7:0] n149;
wire            n150;
wire      [7:0] n151;
wire            n152;
wire      [7:0] n153;
wire            n154;
wire      [7:0] n155;
wire            n156;
wire      [7:0] n157;
wire            n158;
wire      [7:0] n159;
wire      [7:0] n160;
wire      [7:0] n161;
wire      [7:0] n162;
wire      [7:0] n163;
wire      [7:0] n164;
wire      [7:0] n165;
wire      [7:0] n166;
wire      [7:0] n167;
wire      [7:0] n168;
wire      [7:0] n169;
wire      [7:0] n170;
wire      [7:0] n171;
wire      [7:0] n172;
wire      [7:0] n173;
wire      [7:0] n174;
wire      [7:0] n175;
wire      [7:0] n176;
wire      [7:0] n177;
wire      [7:0] n178;
wire      [7:0] n179;
wire      [7:0] n180;
wire      [7:0] n181;
wire      [7:0] n182;
wire      [7:0] n183;
wire      [7:0] n184;
wire      [7:0] n185;
wire      [7:0] n186;
wire      [7:0] n187;
wire      [7:0] n188;
wire      [7:0] n189;
wire      [7:0] n190;
wire      [7:0] n191;
wire      [7:0] n192;
wire      [7:0] n193;
wire      [7:0] n194;
wire      [7:0] n195;
wire      [7:0] n196;
wire      [7:0] n197;
wire      [7:0] n198;
wire      [7:0] n199;
wire      [7:0] n200;
wire      [7:0] n201;
wire      [7:0] n202;
wire      [7:0] n203;
wire      [7:0] n204;
wire      [7:0] n205;
wire      [7:0] n206;
wire      [7:0] n207;
wire      [7:0] n208;
wire      [7:0] n209;
wire      [7:0] n210;
wire      [7:0] n211;
wire      [7:0] n212;
wire      [7:0] n213;
wire      [7:0] n214;
wire      [7:0] n215;
wire      [7:0] n216;
wire     [15:0] n217;
wire     [23:0] n218;
wire     [31:0] n219;
wire     [39:0] n220;
wire     [47:0] n221;
wire     [55:0] n222;
wire     [63:0] n223;
wire     [71:0] n224;
wire     [71:0] n225;
wire     [71:0] n226;
wire     [71:0] n227;
wire     [71:0] n228;
wire     [71:0] n229;
wire     [71:0] n230;
wire     [71:0] n231;
wire     [71:0] n232;
wire     [71:0] n233;
wire     [71:0] n234;
wire     [71:0] n235;
wire            n236;
wire            n237;
wire            n238;
wire            n239;
wire            n240;
wire            n241;
wire            n242;
wire            n243;
wire            n244;
wire            n245;
wire            n246;
wire            n247;
wire            n248;
wire            n249;
wire            n250;
wire            n251;
wire      [7:0] n252;
wire      [7:0] n253;
wire      [7:0] n254;
wire      [7:0] n255;
wire      [7:0] n256;
wire      [7:0] n257;
wire      [7:0] n258;
wire      [7:0] n259;
wire      [7:0] n260;
wire     [15:0] n261;
wire     [23:0] n262;
wire     [31:0] n263;
wire     [39:0] n264;
wire     [47:0] n265;
wire     [55:0] n266;
wire     [63:0] n267;
wire     [71:0] n268;
wire      [7:0] n269;
wire      [7:0] n270;
wire      [7:0] n271;
wire      [7:0] n272;
wire      [7:0] n273;
wire      [7:0] n274;
wire      [7:0] n275;
wire      [7:0] n276;
wire      [7:0] n277;
wire     [15:0] n278;
wire     [23:0] n279;
wire     [31:0] n280;
wire     [39:0] n281;
wire     [47:0] n282;
wire     [55:0] n283;
wire     [63:0] n284;
wire     [71:0] n285;
wire      [7:0] n286;
wire      [7:0] n287;
wire      [7:0] n288;
wire      [7:0] n289;
wire      [7:0] n290;
wire      [7:0] n291;
wire      [7:0] n292;
wire      [7:0] n293;
wire      [7:0] n294;
wire     [15:0] n295;
wire     [23:0] n296;
wire     [31:0] n297;
wire     [39:0] n298;
wire     [47:0] n299;
wire     [55:0] n300;
wire     [63:0] n301;
wire     [71:0] n302;
wire      [7:0] n303;
wire      [7:0] n304;
wire      [7:0] n305;
wire      [7:0] n306;
wire      [7:0] n307;
wire      [7:0] n308;
wire      [7:0] n309;
wire      [7:0] n310;
wire      [7:0] n311;
wire     [15:0] n312;
wire     [23:0] n313;
wire     [31:0] n314;
wire     [39:0] n315;
wire     [47:0] n316;
wire     [55:0] n317;
wire     [63:0] n318;
wire     [71:0] n319;
wire      [7:0] n320;
wire      [7:0] n321;
wire      [7:0] n322;
wire      [7:0] n323;
wire      [7:0] n324;
wire      [7:0] n325;
wire      [7:0] n326;
wire      [7:0] n327;
wire      [7:0] n328;
wire     [15:0] n329;
wire     [23:0] n330;
wire     [31:0] n331;
wire     [39:0] n332;
wire     [47:0] n333;
wire     [55:0] n334;
wire     [63:0] n335;
wire     [71:0] n336;
wire      [7:0] n337;
wire      [7:0] n338;
wire      [7:0] n339;
wire      [7:0] n340;
wire      [7:0] n341;
wire      [7:0] n342;
wire      [7:0] n343;
wire      [7:0] n344;
wire      [7:0] n345;
wire     [15:0] n346;
wire     [23:0] n347;
wire     [31:0] n348;
wire     [39:0] n349;
wire     [47:0] n350;
wire     [55:0] n351;
wire     [63:0] n352;
wire     [71:0] n353;
wire      [7:0] n354;
wire      [7:0] n355;
wire      [7:0] n356;
wire      [7:0] n357;
wire      [7:0] n358;
wire      [7:0] n359;
wire      [7:0] n360;
wire      [7:0] n361;
wire      [7:0] n362;
wire     [15:0] n363;
wire     [23:0] n364;
wire     [31:0] n365;
wire     [39:0] n366;
wire     [47:0] n367;
wire     [55:0] n368;
wire     [63:0] n369;
wire     [71:0] n370;
wire      [7:0] n371;
wire      [7:0] n372;
wire      [7:0] n373;
wire      [7:0] n374;
wire      [7:0] n375;
wire      [7:0] n376;
wire      [7:0] n377;
wire      [7:0] n378;
wire      [7:0] n379;
wire     [15:0] n380;
wire     [23:0] n381;
wire     [31:0] n382;
wire     [39:0] n383;
wire     [47:0] n384;
wire     [55:0] n385;
wire     [63:0] n386;
wire     [71:0] n387;
wire      [7:0] n388;
wire      [7:0] n389;
wire      [7:0] n390;
wire      [7:0] n391;
wire      [7:0] n392;
wire      [7:0] n393;
wire      [7:0] n394;
wire      [7:0] n395;
wire      [7:0] n396;
wire     [15:0] n397;
wire     [23:0] n398;
wire     [31:0] n399;
wire     [39:0] n400;
wire     [47:0] n401;
wire     [55:0] n402;
wire     [63:0] n403;
wire     [71:0] n404;
wire    [143:0] n405;
wire    [215:0] n406;
wire    [287:0] n407;
wire    [359:0] n408;
wire    [431:0] n409;
wire    [503:0] n410;
wire    [575:0] n411;
wire    [647:0] n412;
wire    [647:0] n413;
wire    [647:0] n414;
wire    [647:0] n415;
wire    [647:0] n416;
wire    [647:0] n417;
wire    [647:0] n418;
wire    [647:0] n419;
wire    [647:0] n420;
wire    [647:0] n421;
wire    [647:0] n422;
wire    [647:0] n423;
wire            n424;
wire            n425;
wire            n426;
wire            n427;
wire            n428;
wire            n429;
wire            n430;
wire            n431;
wire            n432;
wire            n433;
wire            n434;
wire            n435;
wire      [8:0] LB2D_proc_0_addr0;
wire      [7:0] LB2D_proc_0_data0;
wire            n436;
wire            n437;
wire            n438;
wire            n439;
wire            n440;
wire            n441;
wire            n442;
wire            n443;
wire            n444;
wire            n445;
wire            n446;
wire            n447;
wire            n448;
wire            n449;
wire            n450;
wire            n451;
wire      [8:0] LB2D_proc_1_addr0;
wire      [7:0] LB2D_proc_1_data0;
wire            n452;
wire            n453;
wire            n454;
wire      [8:0] LB2D_proc_2_addr0;
wire      [7:0] LB2D_proc_2_data0;
wire            n455;
wire            n456;
wire            n457;
wire      [8:0] LB2D_proc_3_addr0;
wire      [7:0] LB2D_proc_3_data0;
wire            n458;
wire            n459;
wire            n460;
wire      [8:0] LB2D_proc_4_addr0;
wire      [7:0] LB2D_proc_4_data0;
wire            n461;
wire            n462;
wire            n463;
wire      [8:0] LB2D_proc_5_addr0;
wire      [7:0] LB2D_proc_5_data0;
wire            n464;
wire            n465;
wire            n466;
wire      [8:0] LB2D_proc_6_addr0;
wire      [7:0] LB2D_proc_6_data0;
wire            n467;
wire            n468;
wire            n469;
wire      [8:0] LB2D_proc_7_addr0;
wire      [7:0] LB2D_proc_7_data0;
wire            n470;
wire            n471;
wire            n472;
wire            n473;
reg      [7:0] LB2D_proc_0[511:0];
reg      [7:0] LB2D_proc_1[511:0];
reg      [7:0] LB2D_proc_2[511:0];
reg      [7:0] LB2D_proc_3[511:0];
reg      [7:0] LB2D_proc_4[511:0];
reg      [7:0] LB2D_proc_5[511:0];
reg      [7:0] LB2D_proc_6[511:0];
reg      [7:0] LB2D_proc_7[511:0];
wire clk;
wire rst;
wire step;
assign n0 =  ( slice_stream_empty ) == ( 1'd0 )  ;
assign n1 =  ( stencil_stream_full ) == ( 1'd0 )  ;
assign n2 =  ( n0 ) & ( n1 )  ;
assign n3 =  ( in_stream_empty ) == ( 1'd0 )  ;
assign n4 =  ( slice_stream_full ) == ( 1'd0 )  ;
assign n5 =  ( n3 ) & ( n4 )  ;
assign n6 =  ( arg_1_TREADY ) == ( 1'd0 )  ;
assign n7 =  ( in_stream_full ) == ( 1'd0 )  ;
assign n8 =  ( n6 ) & ( n7 )  ;
assign n9 =  ( arg_0_TREADY ) == ( 1'd1 )  ;
assign n10 =  ( arg_0_TVALID ) == ( 1'd1 )  ;
assign n11 =  ( n9 ) & ( n10 )  ;
assign n12 =  ( arg_1_TVALID ) == ( 1'd0 )  ;
assign n13 =  ( n11 ) & ( n12 )  ;
assign n14 =  ( arg_1_TREADY ) == ( 1'd1 )  ;
assign n15 =  ( arg_1_TVALID ) == ( 1'd1 )  ;
assign n16 =  ( n14 ) & ( n15 )  ;
assign n17 =  ( arg_0_TREADY ) == ( 1'd0 )  ;
assign n18 =  ( n16 ) & ( n17 )  ;
assign n19 =  ( n18 ) ? ( arg_1_TDATA ) : ( LB1D_buff ) ;
assign n20 =  ( n13 ) ? ( arg_1_TDATA ) : ( n19 ) ;
assign n21 =  ( n8 ) ? ( LB1D_buff ) : ( n20 ) ;
assign n22 =  ( n5 ) ? ( LB1D_buff ) : ( n21 ) ;
assign n23 =  ( n2 ) ? ( LB1D_buff ) : ( n22 ) ;
assign n24 =  ( LB2D_proc_w ) < ( 64'd7 )  ;
assign n25 =  ( LB2D_proc_x ) < ( 9'd487 )  ;
assign n26 =  ( LB2D_proc_w ) + ( 64'd1 )  ;
assign n27 =  ( n25 ) ? ( LB2D_proc_w ) : ( n26 ) ;
assign n28 =  ( n24 ) ? ( n27 ) : ( 64'd0 ) ;
assign n29 =  ( n18 ) ? ( LB2D_proc_w ) : ( LB2D_proc_w ) ;
assign n30 =  ( n13 ) ? ( LB2D_proc_w ) : ( n29 ) ;
assign n31 =  ( n8 ) ? ( LB2D_proc_w ) : ( n30 ) ;
assign n32 =  ( n5 ) ? ( n28 ) : ( n31 ) ;
assign n33 =  ( n2 ) ? ( LB2D_proc_w ) : ( n32 ) ;
assign n34 =  ( LB2D_proc_x ) + ( 9'd1 )  ;
assign n35 =  ( n25 ) ? ( n34 ) : ( 9'd0 ) ;
assign n36 =  ( n18 ) ? ( LB2D_proc_x ) : ( LB2D_proc_x ) ;
assign n37 =  ( n13 ) ? ( LB2D_proc_x ) : ( n36 ) ;
assign n38 =  ( n8 ) ? ( LB2D_proc_x ) : ( n37 ) ;
assign n39 =  ( n5 ) ? ( n35 ) : ( n38 ) ;
assign n40 =  ( n2 ) ? ( LB2D_proc_x ) : ( n39 ) ;
assign n41 =  ( LB2D_proc_y ) < ( 10'd487 )  ;
assign n42 =  ( LB2D_proc_y ) + ( 10'd1 )  ;
assign n43 =  ( n25 ) ? ( LB2D_proc_y ) : ( n42 ) ;
assign n44 =  ( n41 ) ? ( n43 ) : ( 10'd487 ) ;
assign n45 =  ( n18 ) ? ( LB2D_proc_y ) : ( LB2D_proc_y ) ;
assign n46 =  ( n13 ) ? ( LB2D_proc_y ) : ( n45 ) ;
assign n47 =  ( n8 ) ? ( LB2D_proc_y ) : ( n46 ) ;
assign n48 =  ( n5 ) ? ( n44 ) : ( n47 ) ;
assign n49 =  ( n2 ) ? ( LB2D_proc_y ) : ( n48 ) ;
assign n50 =  ( slice_stream_full ) == ( 1'd1 )  ;
assign n51 =  ( n50 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n52 =  ( n18 ) ? ( LB2D_shift_0 ) : ( LB2D_shift_0 ) ;
assign n53 =  ( n13 ) ? ( LB2D_shift_0 ) : ( n52 ) ;
assign n54 =  ( n8 ) ? ( LB2D_shift_0 ) : ( n53 ) ;
assign n55 =  ( n5 ) ? ( LB2D_shift_0 ) : ( n54 ) ;
assign n56 =  ( n2 ) ? ( n51 ) : ( n55 ) ;
assign n57 =  ( n18 ) ? ( LB2D_shift_1 ) : ( LB2D_shift_1 ) ;
assign n58 =  ( n13 ) ? ( LB2D_shift_1 ) : ( n57 ) ;
assign n59 =  ( n8 ) ? ( LB2D_shift_1 ) : ( n58 ) ;
assign n60 =  ( n5 ) ? ( LB2D_shift_1 ) : ( n59 ) ;
assign n61 =  ( n2 ) ? ( LB2D_shift_0 ) : ( n60 ) ;
assign n62 =  ( n18 ) ? ( LB2D_shift_2 ) : ( LB2D_shift_2 ) ;
assign n63 =  ( n13 ) ? ( LB2D_shift_2 ) : ( n62 ) ;
assign n64 =  ( n8 ) ? ( LB2D_shift_2 ) : ( n63 ) ;
assign n65 =  ( n5 ) ? ( LB2D_shift_2 ) : ( n64 ) ;
assign n66 =  ( n2 ) ? ( LB2D_shift_1 ) : ( n65 ) ;
assign n67 =  ( n18 ) ? ( LB2D_shift_3 ) : ( LB2D_shift_3 ) ;
assign n68 =  ( n13 ) ? ( LB2D_shift_3 ) : ( n67 ) ;
assign n69 =  ( n8 ) ? ( LB2D_shift_3 ) : ( n68 ) ;
assign n70 =  ( n5 ) ? ( LB2D_shift_3 ) : ( n69 ) ;
assign n71 =  ( n2 ) ? ( LB2D_shift_2 ) : ( n70 ) ;
assign n72 =  ( n18 ) ? ( LB2D_shift_4 ) : ( LB2D_shift_4 ) ;
assign n73 =  ( n13 ) ? ( LB2D_shift_4 ) : ( n72 ) ;
assign n74 =  ( n8 ) ? ( LB2D_shift_4 ) : ( n73 ) ;
assign n75 =  ( n5 ) ? ( LB2D_shift_4 ) : ( n74 ) ;
assign n76 =  ( n2 ) ? ( LB2D_shift_3 ) : ( n75 ) ;
assign n77 =  ( n18 ) ? ( LB2D_shift_5 ) : ( LB2D_shift_5 ) ;
assign n78 =  ( n13 ) ? ( LB2D_shift_5 ) : ( n77 ) ;
assign n79 =  ( n8 ) ? ( LB2D_shift_5 ) : ( n78 ) ;
assign n80 =  ( n5 ) ? ( LB2D_shift_5 ) : ( n79 ) ;
assign n81 =  ( n2 ) ? ( LB2D_shift_4 ) : ( n80 ) ;
assign n82 =  ( n18 ) ? ( LB2D_shift_6 ) : ( LB2D_shift_6 ) ;
assign n83 =  ( n13 ) ? ( LB2D_shift_6 ) : ( n82 ) ;
assign n84 =  ( n8 ) ? ( LB2D_shift_6 ) : ( n83 ) ;
assign n85 =  ( n5 ) ? ( LB2D_shift_6 ) : ( n84 ) ;
assign n86 =  ( n2 ) ? ( LB2D_shift_5 ) : ( n85 ) ;
assign n87 =  ( n18 ) ? ( LB2D_shift_7 ) : ( LB2D_shift_7 ) ;
assign n88 =  ( n13 ) ? ( LB2D_shift_7 ) : ( n87 ) ;
assign n89 =  ( n8 ) ? ( LB2D_shift_7 ) : ( n88 ) ;
assign n90 =  ( n5 ) ? ( LB2D_shift_7 ) : ( n89 ) ;
assign n91 =  ( n2 ) ? ( LB2D_shift_6 ) : ( n90 ) ;
assign n92 =  ( LB2D_shift_x ) < ( 9'd487 )  ;
assign n93 =  ( LB2D_shift_x ) + ( 9'd1 )  ;
assign n94 =  ( n92 ) ? ( n93 ) : ( 9'd0 ) ;
assign n95 =  ( n18 ) ? ( LB2D_shift_x ) : ( LB2D_shift_x ) ;
assign n96 =  ( n13 ) ? ( LB2D_shift_x ) : ( n95 ) ;
assign n97 =  ( n8 ) ? ( LB2D_shift_x ) : ( n96 ) ;
assign n98 =  ( n5 ) ? ( LB2D_shift_x ) : ( n97 ) ;
assign n99 =  ( n2 ) ? ( n94 ) : ( n98 ) ;
assign n100 =  ( n18 ) ? ( LB2D_shift_y ) : ( LB2D_shift_y ) ;
assign n101 =  ( n13 ) ? ( LB2D_shift_y ) : ( n100 ) ;
assign n102 =  ( n8 ) ? ( LB2D_shift_y ) : ( n101 ) ;
assign n103 =  ( n5 ) ? ( LB2D_shift_y ) : ( n102 ) ;
assign n104 =  ( n2 ) ? ( LB2D_shift_y ) : ( n103 ) ;
assign n105 =  ( n18 ) ? ( arg_0_TDATA ) : ( arg_0_TDATA ) ;
assign n106 =  ( n13 ) ? ( arg_0_TDATA ) : ( n105 ) ;
assign n107 =  ( n8 ) ? ( arg_0_TDATA ) : ( n106 ) ;
assign n108 =  ( n5 ) ? ( arg_0_TDATA ) : ( n107 ) ;
assign n109 =  ( n2 ) ? ( arg_0_TDATA ) : ( n108 ) ;
assign n110 =  ( n18 ) ? ( arg_0_TVALID ) : ( arg_0_TVALID ) ;
assign n111 =  ( n13 ) ? ( 1'd0 ) : ( n110 ) ;
assign n112 =  ( n8 ) ? ( arg_0_TVALID ) : ( n111 ) ;
assign n113 =  ( n5 ) ? ( arg_0_TVALID ) : ( n112 ) ;
assign n114 =  ( n2 ) ? ( arg_0_TVALID ) : ( n113 ) ;
assign n115 =  ( n18 ) ? ( 1'd0 ) : ( arg_1_TREADY ) ;
assign n116 =  ( n13 ) ? ( 1'd0 ) : ( n115 ) ;
assign n117 =  ( n8 ) ? ( 1'd1 ) : ( n116 ) ;
assign n118 =  ( n5 ) ? ( arg_1_TREADY ) : ( n117 ) ;
assign n119 =  ( n2 ) ? ( arg_1_TREADY ) : ( n118 ) ;
assign n120 =  ( n18 ) ? ( in_stream_buff_0 ) : ( in_stream_buff_0 ) ;
assign n121 =  ( n13 ) ? ( in_stream_buff_0 ) : ( n120 ) ;
assign n122 =  ( n8 ) ? ( LB1D_buff ) : ( n121 ) ;
assign n123 =  ( n5 ) ? ( in_stream_buff_0 ) : ( n122 ) ;
assign n124 =  ( n2 ) ? ( in_stream_buff_0 ) : ( n123 ) ;
assign n125 =  ( n18 ) ? ( in_stream_buff_1 ) : ( in_stream_buff_1 ) ;
assign n126 =  ( n13 ) ? ( in_stream_buff_1 ) : ( n125 ) ;
assign n127 =  ( n8 ) ? ( in_stream_buff_0 ) : ( n126 ) ;
assign n128 =  ( n5 ) ? ( in_stream_buff_1 ) : ( n127 ) ;
assign n129 =  ( n2 ) ? ( in_stream_buff_1 ) : ( n128 ) ;
assign n130 =  ( in_stream_full ) == ( 1'd1 )  ;
assign n131 =  ( n130 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n132 =  ( n18 ) ? ( in_stream_empty ) : ( in_stream_empty ) ;
assign n133 =  ( n13 ) ? ( in_stream_empty ) : ( n132 ) ;
assign n134 =  ( n8 ) ? ( 1'd0 ) : ( n133 ) ;
assign n135 =  ( n5 ) ? ( n131 ) : ( n134 ) ;
assign n136 =  ( n2 ) ? ( in_stream_empty ) : ( n135 ) ;
assign n137 =  ( in_stream_empty ) == ( 1'd1 )  ;
assign n138 =  ( n137 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n139 =  ( n18 ) ? ( in_stream_full ) : ( in_stream_full ) ;
assign n140 =  ( n13 ) ? ( in_stream_full ) : ( n139 ) ;
assign n141 =  ( n8 ) ? ( n138 ) : ( n140 ) ;
assign n142 =  ( n5 ) ? ( 1'd0 ) : ( n141 ) ;
assign n143 =  ( n2 ) ? ( in_stream_full ) : ( n142 ) ;
assign n144 =  ( LB2D_proc_y ) >= ( 10'd8 )  ;
assign n145 =  ( n130 ) ? ( in_stream_buff_1 ) : ( in_stream_buff_0 ) ;
assign n146 =  ( LB2D_proc_w ) == ( 64'd0 )  ;
assign n147 =  (  LB2D_proc_7 [ LB2D_proc_x ] )  ;
assign n148 =  ( LB2D_proc_w ) == ( 64'd1 )  ;
assign n149 =  (  LB2D_proc_0 [ LB2D_proc_x ] )  ;
assign n150 =  ( LB2D_proc_w ) == ( 64'd2 )  ;
assign n151 =  (  LB2D_proc_1 [ LB2D_proc_x ] )  ;
assign n152 =  ( LB2D_proc_w ) == ( 64'd3 )  ;
assign n153 =  (  LB2D_proc_2 [ LB2D_proc_x ] )  ;
assign n154 =  ( LB2D_proc_w ) == ( 64'd4 )  ;
assign n155 =  (  LB2D_proc_3 [ LB2D_proc_x ] )  ;
assign n156 =  ( LB2D_proc_w ) == ( 64'd5 )  ;
assign n157 =  (  LB2D_proc_4 [ LB2D_proc_x ] )  ;
assign n158 =  ( LB2D_proc_w ) == ( 64'd6 )  ;
assign n159 =  (  LB2D_proc_5 [ LB2D_proc_x ] )  ;
assign n160 =  (  LB2D_proc_6 [ LB2D_proc_x ] )  ;
assign n161 =  ( n158 ) ? ( n159 ) : ( n160 ) ;
assign n162 =  ( n156 ) ? ( n157 ) : ( n161 ) ;
assign n163 =  ( n154 ) ? ( n155 ) : ( n162 ) ;
assign n164 =  ( n152 ) ? ( n153 ) : ( n163 ) ;
assign n165 =  ( n150 ) ? ( n151 ) : ( n164 ) ;
assign n166 =  ( n148 ) ? ( n149 ) : ( n165 ) ;
assign n167 =  ( n146 ) ? ( n147 ) : ( n166 ) ;
assign n168 =  ( n158 ) ? ( n157 ) : ( n159 ) ;
assign n169 =  ( n156 ) ? ( n155 ) : ( n168 ) ;
assign n170 =  ( n154 ) ? ( n153 ) : ( n169 ) ;
assign n171 =  ( n152 ) ? ( n151 ) : ( n170 ) ;
assign n172 =  ( n150 ) ? ( n149 ) : ( n171 ) ;
assign n173 =  ( n148 ) ? ( n147 ) : ( n172 ) ;
assign n174 =  ( n146 ) ? ( n160 ) : ( n173 ) ;
assign n175 =  ( n158 ) ? ( n155 ) : ( n157 ) ;
assign n176 =  ( n156 ) ? ( n153 ) : ( n175 ) ;
assign n177 =  ( n154 ) ? ( n151 ) : ( n176 ) ;
assign n178 =  ( n152 ) ? ( n149 ) : ( n177 ) ;
assign n179 =  ( n150 ) ? ( n147 ) : ( n178 ) ;
assign n180 =  ( n148 ) ? ( n160 ) : ( n179 ) ;
assign n181 =  ( n146 ) ? ( n159 ) : ( n180 ) ;
assign n182 =  ( n158 ) ? ( n153 ) : ( n155 ) ;
assign n183 =  ( n156 ) ? ( n151 ) : ( n182 ) ;
assign n184 =  ( n154 ) ? ( n149 ) : ( n183 ) ;
assign n185 =  ( n152 ) ? ( n147 ) : ( n184 ) ;
assign n186 =  ( n150 ) ? ( n160 ) : ( n185 ) ;
assign n187 =  ( n148 ) ? ( n159 ) : ( n186 ) ;
assign n188 =  ( n146 ) ? ( n157 ) : ( n187 ) ;
assign n189 =  ( n158 ) ? ( n151 ) : ( n153 ) ;
assign n190 =  ( n156 ) ? ( n149 ) : ( n189 ) ;
assign n191 =  ( n154 ) ? ( n147 ) : ( n190 ) ;
assign n192 =  ( n152 ) ? ( n160 ) : ( n191 ) ;
assign n193 =  ( n150 ) ? ( n159 ) : ( n192 ) ;
assign n194 =  ( n148 ) ? ( n157 ) : ( n193 ) ;
assign n195 =  ( n146 ) ? ( n155 ) : ( n194 ) ;
assign n196 =  ( n158 ) ? ( n149 ) : ( n151 ) ;
assign n197 =  ( n156 ) ? ( n147 ) : ( n196 ) ;
assign n198 =  ( n154 ) ? ( n160 ) : ( n197 ) ;
assign n199 =  ( n152 ) ? ( n159 ) : ( n198 ) ;
assign n200 =  ( n150 ) ? ( n157 ) : ( n199 ) ;
assign n201 =  ( n148 ) ? ( n155 ) : ( n200 ) ;
assign n202 =  ( n146 ) ? ( n153 ) : ( n201 ) ;
assign n203 =  ( n158 ) ? ( n147 ) : ( n149 ) ;
assign n204 =  ( n156 ) ? ( n160 ) : ( n203 ) ;
assign n205 =  ( n154 ) ? ( n159 ) : ( n204 ) ;
assign n206 =  ( n152 ) ? ( n157 ) : ( n205 ) ;
assign n207 =  ( n150 ) ? ( n155 ) : ( n206 ) ;
assign n208 =  ( n148 ) ? ( n153 ) : ( n207 ) ;
assign n209 =  ( n146 ) ? ( n151 ) : ( n208 ) ;
assign n210 =  ( n158 ) ? ( n160 ) : ( n147 ) ;
assign n211 =  ( n156 ) ? ( n159 ) : ( n210 ) ;
assign n212 =  ( n154 ) ? ( n157 ) : ( n211 ) ;
assign n213 =  ( n152 ) ? ( n155 ) : ( n212 ) ;
assign n214 =  ( n150 ) ? ( n153 ) : ( n213 ) ;
assign n215 =  ( n148 ) ? ( n151 ) : ( n214 ) ;
assign n216 =  ( n146 ) ? ( n149 ) : ( n215 ) ;
assign n217 =  { ( n209 ) , ( n216 ) }  ;
assign n218 =  { ( n202 ) , ( n217 ) }  ;
assign n219 =  { ( n195 ) , ( n218 ) }  ;
assign n220 =  { ( n188 ) , ( n219 ) }  ;
assign n221 =  { ( n181 ) , ( n220 ) }  ;
assign n222 =  { ( n174 ) , ( n221 ) }  ;
assign n223 =  { ( n167 ) , ( n222 ) }  ;
assign n224 =  { ( n145 ) , ( n223 ) }  ;
assign n225 =  ( n144 ) ? ( n224 ) : ( slice_stream_buff_0 ) ;
assign n226 =  ( n18 ) ? ( slice_stream_buff_0 ) : ( slice_stream_buff_0 ) ;
assign n227 =  ( n13 ) ? ( slice_stream_buff_0 ) : ( n226 ) ;
assign n228 =  ( n8 ) ? ( slice_stream_buff_0 ) : ( n227 ) ;
assign n229 =  ( n5 ) ? ( n225 ) : ( n228 ) ;
assign n230 =  ( n2 ) ? ( slice_stream_buff_0 ) : ( n229 ) ;
assign n231 =  ( n18 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_1 ) ;
assign n232 =  ( n13 ) ? ( slice_stream_buff_1 ) : ( n231 ) ;
assign n233 =  ( n8 ) ? ( slice_stream_buff_1 ) : ( n232 ) ;
assign n234 =  ( n5 ) ? ( slice_stream_buff_0 ) : ( n233 ) ;
assign n235 =  ( n2 ) ? ( slice_stream_buff_1 ) : ( n234 ) ;
assign n236 =  ( n50 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n237 =  ( n144 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n238 =  ( n18 ) ? ( slice_stream_empty ) : ( slice_stream_empty ) ;
assign n239 =  ( n13 ) ? ( slice_stream_empty ) : ( n238 ) ;
assign n240 =  ( n8 ) ? ( slice_stream_empty ) : ( n239 ) ;
assign n241 =  ( n5 ) ? ( n237 ) : ( n240 ) ;
assign n242 =  ( n2 ) ? ( n236 ) : ( n241 ) ;
assign n243 =  ( slice_stream_empty ) == ( 1'd1 )  ;
assign n244 =  ( n243 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n245 =  ( n144 ) ? ( n244 ) : ( 1'd0 ) ;
assign n246 =  ( n18 ) ? ( slice_stream_full ) : ( slice_stream_full ) ;
assign n247 =  ( n13 ) ? ( slice_stream_full ) : ( n246 ) ;
assign n248 =  ( n8 ) ? ( slice_stream_full ) : ( n247 ) ;
assign n249 =  ( n5 ) ? ( n245 ) : ( n248 ) ;
assign n250 =  ( n2 ) ? ( 1'd0 ) : ( n249 ) ;
assign n251 =  ( LB2D_shift_x ) >= ( 9'd8 )  ;
assign n252 = n51[71:64] ;
assign n253 = LB2D_shift_0[71:64] ;
assign n254 = LB2D_shift_1[71:64] ;
assign n255 = LB2D_shift_2[71:64] ;
assign n256 = LB2D_shift_3[71:64] ;
assign n257 = LB2D_shift_4[71:64] ;
assign n258 = LB2D_shift_5[71:64] ;
assign n259 = LB2D_shift_6[71:64] ;
assign n260 = LB2D_shift_7[71:64] ;
assign n261 =  { ( n259 ) , ( n260 ) }  ;
assign n262 =  { ( n258 ) , ( n261 ) }  ;
assign n263 =  { ( n257 ) , ( n262 ) }  ;
assign n264 =  { ( n256 ) , ( n263 ) }  ;
assign n265 =  { ( n255 ) , ( n264 ) }  ;
assign n266 =  { ( n254 ) , ( n265 ) }  ;
assign n267 =  { ( n253 ) , ( n266 ) }  ;
assign n268 =  { ( n252 ) , ( n267 ) }  ;
assign n269 = n51[63:56] ;
assign n270 = LB2D_shift_0[63:56] ;
assign n271 = LB2D_shift_1[63:56] ;
assign n272 = LB2D_shift_2[63:56] ;
assign n273 = LB2D_shift_3[63:56] ;
assign n274 = LB2D_shift_4[63:56] ;
assign n275 = LB2D_shift_5[63:56] ;
assign n276 = LB2D_shift_6[63:56] ;
assign n277 = LB2D_shift_7[63:56] ;
assign n278 =  { ( n276 ) , ( n277 ) }  ;
assign n279 =  { ( n275 ) , ( n278 ) }  ;
assign n280 =  { ( n274 ) , ( n279 ) }  ;
assign n281 =  { ( n273 ) , ( n280 ) }  ;
assign n282 =  { ( n272 ) , ( n281 ) }  ;
assign n283 =  { ( n271 ) , ( n282 ) }  ;
assign n284 =  { ( n270 ) , ( n283 ) }  ;
assign n285 =  { ( n269 ) , ( n284 ) }  ;
assign n286 = n51[55:48] ;
assign n287 = LB2D_shift_0[55:48] ;
assign n288 = LB2D_shift_1[55:48] ;
assign n289 = LB2D_shift_2[55:48] ;
assign n290 = LB2D_shift_3[55:48] ;
assign n291 = LB2D_shift_4[55:48] ;
assign n292 = LB2D_shift_5[55:48] ;
assign n293 = LB2D_shift_6[55:48] ;
assign n294 = LB2D_shift_7[55:48] ;
assign n295 =  { ( n293 ) , ( n294 ) }  ;
assign n296 =  { ( n292 ) , ( n295 ) }  ;
assign n297 =  { ( n291 ) , ( n296 ) }  ;
assign n298 =  { ( n290 ) , ( n297 ) }  ;
assign n299 =  { ( n289 ) , ( n298 ) }  ;
assign n300 =  { ( n288 ) , ( n299 ) }  ;
assign n301 =  { ( n287 ) , ( n300 ) }  ;
assign n302 =  { ( n286 ) , ( n301 ) }  ;
assign n303 = n51[47:40] ;
assign n304 = LB2D_shift_0[47:40] ;
assign n305 = LB2D_shift_1[47:40] ;
assign n306 = LB2D_shift_2[47:40] ;
assign n307 = LB2D_shift_3[47:40] ;
assign n308 = LB2D_shift_4[47:40] ;
assign n309 = LB2D_shift_5[47:40] ;
assign n310 = LB2D_shift_6[47:40] ;
assign n311 = LB2D_shift_7[47:40] ;
assign n312 =  { ( n310 ) , ( n311 ) }  ;
assign n313 =  { ( n309 ) , ( n312 ) }  ;
assign n314 =  { ( n308 ) , ( n313 ) }  ;
assign n315 =  { ( n307 ) , ( n314 ) }  ;
assign n316 =  { ( n306 ) , ( n315 ) }  ;
assign n317 =  { ( n305 ) , ( n316 ) }  ;
assign n318 =  { ( n304 ) , ( n317 ) }  ;
assign n319 =  { ( n303 ) , ( n318 ) }  ;
assign n320 = n51[39:32] ;
assign n321 = LB2D_shift_0[39:32] ;
assign n322 = LB2D_shift_1[39:32] ;
assign n323 = LB2D_shift_2[39:32] ;
assign n324 = LB2D_shift_3[39:32] ;
assign n325 = LB2D_shift_4[39:32] ;
assign n326 = LB2D_shift_5[39:32] ;
assign n327 = LB2D_shift_6[39:32] ;
assign n328 = LB2D_shift_7[39:32] ;
assign n329 =  { ( n327 ) , ( n328 ) }  ;
assign n330 =  { ( n326 ) , ( n329 ) }  ;
assign n331 =  { ( n325 ) , ( n330 ) }  ;
assign n332 =  { ( n324 ) , ( n331 ) }  ;
assign n333 =  { ( n323 ) , ( n332 ) }  ;
assign n334 =  { ( n322 ) , ( n333 ) }  ;
assign n335 =  { ( n321 ) , ( n334 ) }  ;
assign n336 =  { ( n320 ) , ( n335 ) }  ;
assign n337 = n51[31:24] ;
assign n338 = LB2D_shift_0[31:24] ;
assign n339 = LB2D_shift_1[31:24] ;
assign n340 = LB2D_shift_2[31:24] ;
assign n341 = LB2D_shift_3[31:24] ;
assign n342 = LB2D_shift_4[31:24] ;
assign n343 = LB2D_shift_5[31:24] ;
assign n344 = LB2D_shift_6[31:24] ;
assign n345 = LB2D_shift_7[31:24] ;
assign n346 =  { ( n344 ) , ( n345 ) }  ;
assign n347 =  { ( n343 ) , ( n346 ) }  ;
assign n348 =  { ( n342 ) , ( n347 ) }  ;
assign n349 =  { ( n341 ) , ( n348 ) }  ;
assign n350 =  { ( n340 ) , ( n349 ) }  ;
assign n351 =  { ( n339 ) , ( n350 ) }  ;
assign n352 =  { ( n338 ) , ( n351 ) }  ;
assign n353 =  { ( n337 ) , ( n352 ) }  ;
assign n354 = n51[23:16] ;
assign n355 = LB2D_shift_0[23:16] ;
assign n356 = LB2D_shift_1[23:16] ;
assign n357 = LB2D_shift_2[23:16] ;
assign n358 = LB2D_shift_3[23:16] ;
assign n359 = LB2D_shift_4[23:16] ;
assign n360 = LB2D_shift_5[23:16] ;
assign n361 = LB2D_shift_6[23:16] ;
assign n362 = LB2D_shift_7[23:16] ;
assign n363 =  { ( n361 ) , ( n362 ) }  ;
assign n364 =  { ( n360 ) , ( n363 ) }  ;
assign n365 =  { ( n359 ) , ( n364 ) }  ;
assign n366 =  { ( n358 ) , ( n365 ) }  ;
assign n367 =  { ( n357 ) , ( n366 ) }  ;
assign n368 =  { ( n356 ) , ( n367 ) }  ;
assign n369 =  { ( n355 ) , ( n368 ) }  ;
assign n370 =  { ( n354 ) , ( n369 ) }  ;
assign n371 = n51[15:8] ;
assign n372 = LB2D_shift_0[15:8] ;
assign n373 = LB2D_shift_1[15:8] ;
assign n374 = LB2D_shift_2[15:8] ;
assign n375 = LB2D_shift_3[15:8] ;
assign n376 = LB2D_shift_4[15:8] ;
assign n377 = LB2D_shift_5[15:8] ;
assign n378 = LB2D_shift_6[15:8] ;
assign n379 = LB2D_shift_7[15:8] ;
assign n380 =  { ( n378 ) , ( n379 ) }  ;
assign n381 =  { ( n377 ) , ( n380 ) }  ;
assign n382 =  { ( n376 ) , ( n381 ) }  ;
assign n383 =  { ( n375 ) , ( n382 ) }  ;
assign n384 =  { ( n374 ) , ( n383 ) }  ;
assign n385 =  { ( n373 ) , ( n384 ) }  ;
assign n386 =  { ( n372 ) , ( n385 ) }  ;
assign n387 =  { ( n371 ) , ( n386 ) }  ;
assign n388 = n51[7:0] ;
assign n389 = LB2D_shift_0[7:0] ;
assign n390 = LB2D_shift_1[7:0] ;
assign n391 = LB2D_shift_2[7:0] ;
assign n392 = LB2D_shift_3[7:0] ;
assign n393 = LB2D_shift_4[7:0] ;
assign n394 = LB2D_shift_5[7:0] ;
assign n395 = LB2D_shift_6[7:0] ;
assign n396 = LB2D_shift_7[7:0] ;
assign n397 =  { ( n395 ) , ( n396 ) }  ;
assign n398 =  { ( n394 ) , ( n397 ) }  ;
assign n399 =  { ( n393 ) , ( n398 ) }  ;
assign n400 =  { ( n392 ) , ( n399 ) }  ;
assign n401 =  { ( n391 ) , ( n400 ) }  ;
assign n402 =  { ( n390 ) , ( n401 ) }  ;
assign n403 =  { ( n389 ) , ( n402 ) }  ;
assign n404 =  { ( n388 ) , ( n403 ) }  ;
assign n405 =  { ( n387 ) , ( n404 ) }  ;
assign n406 =  { ( n370 ) , ( n405 ) }  ;
assign n407 =  { ( n353 ) , ( n406 ) }  ;
assign n408 =  { ( n336 ) , ( n407 ) }  ;
assign n409 =  { ( n319 ) , ( n408 ) }  ;
assign n410 =  { ( n302 ) , ( n409 ) }  ;
assign n411 =  { ( n285 ) , ( n410 ) }  ;
assign n412 =  { ( n268 ) , ( n411 ) }  ;
assign n413 =  ( n251 ) ? ( n412 ) : ( stencil_stream_buff_0 ) ;
assign n414 =  ( n18 ) ? ( stencil_stream_buff_0 ) : ( stencil_stream_buff_0 ) ;
assign n415 =  ( n13 ) ? ( stencil_stream_buff_0 ) : ( n414 ) ;
assign n416 =  ( n8 ) ? ( stencil_stream_buff_0 ) : ( n415 ) ;
assign n417 =  ( n5 ) ? ( stencil_stream_buff_0 ) : ( n416 ) ;
assign n418 =  ( n2 ) ? ( n413 ) : ( n417 ) ;
assign n419 =  ( n18 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_1 ) ;
assign n420 =  ( n13 ) ? ( stencil_stream_buff_1 ) : ( n419 ) ;
assign n421 =  ( n8 ) ? ( stencil_stream_buff_1 ) : ( n420 ) ;
assign n422 =  ( n5 ) ? ( stencil_stream_buff_1 ) : ( n421 ) ;
assign n423 =  ( n2 ) ? ( stencil_stream_buff_0 ) : ( n422 ) ;
assign n424 =  ( n18 ) ? ( stencil_stream_empty ) : ( stencil_stream_empty ) ;
assign n425 =  ( n13 ) ? ( stencil_stream_empty ) : ( n424 ) ;
assign n426 =  ( n8 ) ? ( stencil_stream_empty ) : ( n425 ) ;
assign n427 =  ( n5 ) ? ( stencil_stream_empty ) : ( n426 ) ;
assign n428 =  ( stencil_stream_empty ) == ( 1'd1 )  ;
assign n429 =  ( n428 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n430 =  ( n251 ) ? ( n429 ) : ( 1'd0 ) ;
assign n431 =  ( n18 ) ? ( stencil_stream_full ) : ( stencil_stream_full ) ;
assign n432 =  ( n13 ) ? ( stencil_stream_full ) : ( n431 ) ;
assign n433 =  ( n8 ) ? ( stencil_stream_full ) : ( n432 ) ;
assign n434 =  ( n5 ) ? ( stencil_stream_full ) : ( n433 ) ;
assign n435 =  ( n2 ) ? ( n430 ) : ( n434 ) ;
assign n436 = ~ ( n2 ) ;
assign n437 = ~ ( n5 ) ;
assign n438 =  ( n436 ) & ( n437 )  ;
assign n439 = ~ ( n8 ) ;
assign n440 =  ( n438 ) & ( n439 )  ;
assign n441 = ~ ( n13 ) ;
assign n442 =  ( n440 ) & ( n441 )  ;
assign n443 = ~ ( n18 ) ;
assign n444 =  ( n442 ) & ( n443 )  ;
assign n445 =  ( n442 ) & ( n18 )  ;
assign n446 =  ( n440 ) & ( n13 )  ;
assign n447 =  ( n438 ) & ( n8 )  ;
assign n448 =  ( n436 ) & ( n5 )  ;
assign n449 = ~ ( n146 ) ;
assign n450 =  ( n448 ) & ( n449 )  ;
assign n451 =  ( n448 ) & ( n146 )  ;
assign LB2D_proc_0_addr0 = n451 ? (LB2D_proc_x) : (0);
assign LB2D_proc_0_data0 = n451 ? (n145) : (LB2D_proc_0[0]);
assign n452 = ~ ( n148 ) ;
assign n453 =  ( n448 ) & ( n452 )  ;
assign n454 =  ( n448 ) & ( n148 )  ;
assign LB2D_proc_1_addr0 = n454 ? (LB2D_proc_x) : (0);
assign LB2D_proc_1_data0 = n454 ? (n145) : (LB2D_proc_1[0]);
assign n455 = ~ ( n150 ) ;
assign n456 =  ( n448 ) & ( n455 )  ;
assign n457 =  ( n448 ) & ( n150 )  ;
assign LB2D_proc_2_addr0 = n457 ? (LB2D_proc_x) : (0);
assign LB2D_proc_2_data0 = n457 ? (n145) : (LB2D_proc_2[0]);
assign n458 = ~ ( n152 ) ;
assign n459 =  ( n448 ) & ( n458 )  ;
assign n460 =  ( n448 ) & ( n152 )  ;
assign LB2D_proc_3_addr0 = n460 ? (LB2D_proc_x) : (0);
assign LB2D_proc_3_data0 = n460 ? (n145) : (LB2D_proc_3[0]);
assign n461 = ~ ( n154 ) ;
assign n462 =  ( n448 ) & ( n461 )  ;
assign n463 =  ( n448 ) & ( n154 )  ;
assign LB2D_proc_4_addr0 = n463 ? (LB2D_proc_x) : (0);
assign LB2D_proc_4_data0 = n463 ? (n145) : (LB2D_proc_4[0]);
assign n464 = ~ ( n156 ) ;
assign n465 =  ( n448 ) & ( n464 )  ;
assign n466 =  ( n448 ) & ( n156 )  ;
assign LB2D_proc_5_addr0 = n466 ? (LB2D_proc_x) : (0);
assign LB2D_proc_5_data0 = n466 ? (n145) : (LB2D_proc_5[0]);
assign n467 = ~ ( n158 ) ;
assign n468 =  ( n448 ) & ( n467 )  ;
assign n469 =  ( n448 ) & ( n158 )  ;
assign LB2D_proc_6_addr0 = n469 ? (LB2D_proc_x) : (0);
assign LB2D_proc_6_data0 = n469 ? (n145) : (LB2D_proc_6[0]);
assign n470 =  ( LB2D_proc_w ) == ( 64'd7 )  ;
assign n471 = ~ ( n470 ) ;
assign n472 =  ( n448 ) & ( n471 )  ;
assign n473 =  ( n448 ) & ( n470 )  ;
assign LB2D_proc_7_addr0 = n473 ? (LB2D_proc_x) : (0);
assign LB2D_proc_7_data0 = n473 ? (n145) : (LB2D_proc_7[0]);
always @(posedge clk) begin
   if(rst) begin
       LB1D_buff <= LB1D_buff;
       LB2D_proc_w <= LB2D_proc_w;
       LB2D_proc_x <= LB2D_proc_x;
       LB2D_proc_y <= LB2D_proc_y;
       LB2D_shift_0 <= LB2D_shift_0;
       LB2D_shift_1 <= LB2D_shift_1;
       LB2D_shift_2 <= LB2D_shift_2;
       LB2D_shift_3 <= LB2D_shift_3;
       LB2D_shift_4 <= LB2D_shift_4;
       LB2D_shift_5 <= LB2D_shift_5;
       LB2D_shift_6 <= LB2D_shift_6;
       LB2D_shift_7 <= LB2D_shift_7;
       LB2D_shift_x <= LB2D_shift_x;
       LB2D_shift_y <= LB2D_shift_y;
       arg_0_TDATA <= arg_0_TDATA;
       arg_0_TVALID <= arg_0_TVALID;
       arg_1_TREADY <= arg_1_TREADY;
       in_stream_buff_0 <= in_stream_buff_0;
       in_stream_buff_1 <= in_stream_buff_1;
       in_stream_empty <= in_stream_empty;
       in_stream_full <= in_stream_full;
       slice_stream_buff_0 <= slice_stream_buff_0;
       slice_stream_buff_1 <= slice_stream_buff_1;
       slice_stream_empty <= slice_stream_empty;
       slice_stream_full <= slice_stream_full;
       stencil_stream_buff_0 <= stencil_stream_buff_0;
       stencil_stream_buff_1 <= stencil_stream_buff_1;
       stencil_stream_empty <= stencil_stream_empty;
       stencil_stream_full <= stencil_stream_full;
   end
   else if(step) begin
       LB1D_buff <= n23;
       LB2D_proc_w <= n33;
       LB2D_proc_x <= n40;
       LB2D_proc_y <= n49;
       LB2D_shift_0 <= n56;
       LB2D_shift_1 <= n61;
       LB2D_shift_2 <= n66;
       LB2D_shift_3 <= n71;
       LB2D_shift_4 <= n76;
       LB2D_shift_5 <= n81;
       LB2D_shift_6 <= n86;
       LB2D_shift_7 <= n91;
       LB2D_shift_x <= n99;
       LB2D_shift_y <= n104;
       arg_0_TDATA <= n109;
       arg_0_TVALID <= n114;
       arg_1_TREADY <= n119;
       in_stream_buff_0 <= n124;
       in_stream_buff_1 <= n129;
       in_stream_empty <= n136;
       in_stream_full <= n143;
       slice_stream_buff_0 <= n230;
       slice_stream_buff_1 <= n235;
       slice_stream_empty <= n242;
       slice_stream_full <= n250;
       stencil_stream_buff_0 <= n418;
       stencil_stream_buff_1 <= n423;
       stencil_stream_empty <= n427;
       stencil_stream_full <= n435;
       LB2D_proc_0 [ LB2D_proc_0_addr0 ] <= LB2D_proc_0_data0;
       LB2D_proc_1 [ LB2D_proc_1_addr0 ] <= LB2D_proc_1_data0;
       LB2D_proc_2 [ LB2D_proc_2_addr0 ] <= LB2D_proc_2_data0;
       LB2D_proc_3 [ LB2D_proc_3_addr0 ] <= LB2D_proc_3_data0;
       LB2D_proc_4 [ LB2D_proc_4_addr0 ] <= LB2D_proc_4_data0;
       LB2D_proc_5 [ LB2D_proc_5_addr0 ] <= LB2D_proc_5_data0;
       LB2D_proc_6 [ LB2D_proc_6_addr0 ] <= LB2D_proc_6_data0;
       LB2D_proc_7 [ LB2D_proc_7_addr0 ] <= LB2D_proc_7_data0;
   end
end
endmodule
