module GB(
arg_0_TREADY,
arg_1_TDATA,
arg_1_TVALID,
LB1D_buff,
LB1D_p_cnt,
LB2D_proc_w,
LB2D_proc_x,
LB2D_proc_y,
LB2D_shift_0,
LB2D_shift_1,
LB2D_shift_2,
LB2D_shift_3,
LB2D_shift_4,
LB2D_shift_5,
LB2D_shift_6,
LB2D_shift_7,
LB2D_shift_x,
LB2D_shift_y,
arg_0_TDATA,
arg_0_TVALID,
arg_1_TREADY,
gb_exit_it_1,
gb_exit_it_2,
gb_exit_it_3,
gb_exit_it_4,
gb_exit_it_5,
gb_exit_it_6,
gb_exit_it_7,
gb_exit_it_8,
gb_p_cnt,
gb_pp_it_1,
gb_pp_it_2,
gb_pp_it_3,
gb_pp_it_4,
gb_pp_it_5,
gb_pp_it_6,
gb_pp_it_7,
gb_pp_it_8,
gb_pp_it_9,
in_stream_buff_0,
in_stream_buff_1,
in_stream_empty,
in_stream_full,
slice_stream_buff_0,
slice_stream_buff_1,
slice_stream_empty,
slice_stream_full,
stencil_stream_buff_0,
stencil_stream_buff_1,
stencil_stream_empty,
stencil_stream_full,
clk,rst,
step
);
input            arg_0_TREADY;
input      [7:0] arg_1_TDATA;
input            arg_1_TVALID;
input clk;
input rst;
input step;
output      [7:0] LB1D_buff;
output     [18:0] LB1D_p_cnt;
output     [63:0] LB2D_proc_w;
output      [8:0] LB2D_proc_x;
output      [9:0] LB2D_proc_y;
output     [71:0] LB2D_shift_0;
output     [71:0] LB2D_shift_1;
output     [71:0] LB2D_shift_2;
output     [71:0] LB2D_shift_3;
output     [71:0] LB2D_shift_4;
output     [71:0] LB2D_shift_5;
output     [71:0] LB2D_shift_6;
output     [71:0] LB2D_shift_7;
output      [8:0] LB2D_shift_x;
output      [9:0] LB2D_shift_y;
output      [7:0] arg_0_TDATA;
output            arg_0_TVALID;
output            arg_1_TREADY;
output            gb_exit_it_1;
output            gb_exit_it_2;
output            gb_exit_it_3;
output            gb_exit_it_4;
output            gb_exit_it_5;
output            gb_exit_it_6;
output            gb_exit_it_7;
output            gb_exit_it_8;
output     [18:0] gb_p_cnt;
output            gb_pp_it_1;
output            gb_pp_it_2;
output            gb_pp_it_3;
output            gb_pp_it_4;
output            gb_pp_it_5;
output            gb_pp_it_6;
output            gb_pp_it_7;
output            gb_pp_it_8;
output            gb_pp_it_9;
output      [7:0] in_stream_buff_0;
output      [7:0] in_stream_buff_1;
output            in_stream_empty;
output            in_stream_full;
output     [71:0] slice_stream_buff_0;
output     [71:0] slice_stream_buff_1;
output            slice_stream_empty;
output            slice_stream_full;
output    [647:0] stencil_stream_buff_0;
output    [647:0] stencil_stream_buff_1;
output            stencil_stream_empty;
output            stencil_stream_full;
reg      [7:0] LB1D_buff;
reg     [18:0] LB1D_p_cnt;
reg     [63:0] LB2D_proc_w;
reg      [8:0] LB2D_proc_x;
reg      [9:0] LB2D_proc_y;
reg     [71:0] LB2D_shift_0;
reg     [71:0] LB2D_shift_1;
reg     [71:0] LB2D_shift_2;
reg     [71:0] LB2D_shift_3;
reg     [71:0] LB2D_shift_4;
reg     [71:0] LB2D_shift_5;
reg     [71:0] LB2D_shift_6;
reg     [71:0] LB2D_shift_7;
reg      [8:0] LB2D_shift_x;
reg      [9:0] LB2D_shift_y;
reg      [7:0] arg_0_TDATA;
reg            arg_0_TVALID;
reg            arg_1_TREADY;
reg            gb_exit_it_1;
reg            gb_exit_it_2;
reg            gb_exit_it_3;
reg            gb_exit_it_4;
reg            gb_exit_it_5;
reg            gb_exit_it_6;
reg            gb_exit_it_7;
reg            gb_exit_it_8;
reg     [18:0] gb_p_cnt;
reg            gb_pp_it_1;
reg            gb_pp_it_2;
reg            gb_pp_it_3;
reg            gb_pp_it_4;
reg            gb_pp_it_5;
reg            gb_pp_it_6;
reg            gb_pp_it_7;
reg            gb_pp_it_8;
reg            gb_pp_it_9;
reg      [7:0] in_stream_buff_0;
reg      [7:0] in_stream_buff_1;
reg            in_stream_empty;
reg            in_stream_full;
reg     [71:0] slice_stream_buff_0;
reg     [71:0] slice_stream_buff_1;
reg            slice_stream_empty;
reg            slice_stream_full;
reg    [647:0] stencil_stream_buff_0;
reg    [647:0] stencil_stream_buff_1;
reg            stencil_stream_empty;
reg            stencil_stream_full;
wire            arg_0_TREADY;
wire      [7:0] arg_1_TDATA;
wire            arg_1_TVALID;
wire            n0;
wire            n1;
wire            n2;
wire            n3;
wire            n4;
wire            n5;
wire            n6;
wire            n7;
wire            n8;
wire            n9;
wire            n10;
wire            n11;
wire            n12;
wire            n13;
wire            n14;
wire            n15;
wire            n16;
wire            n17;
wire            n18;
wire            n19;
wire            n20;
wire            n21;
wire            n22;
wire            n23;
wire            n24;
wire            n25;
wire            n26;
wire            n27;
wire            n28;
wire            n29;
wire            n30;
wire            n31;
wire            n32;
wire            n33;
wire      [7:0] n34;
wire      [7:0] n35;
wire      [7:0] n36;
wire      [7:0] n37;
wire      [7:0] n38;
wire      [7:0] n39;
wire     [18:0] n40;
wire     [18:0] n41;
wire            n42;
wire            n43;
wire     [63:0] n44;
wire     [63:0] n45;
wire     [63:0] n46;
wire     [63:0] n47;
wire     [63:0] n48;
wire     [63:0] n49;
wire     [63:0] n50;
wire     [63:0] n51;
wire     [63:0] n52;
wire      [8:0] n53;
wire      [8:0] n54;
wire      [8:0] n55;
wire      [8:0] n56;
wire      [8:0] n57;
wire      [8:0] n58;
wire      [8:0] n59;
wire      [8:0] n60;
wire            n61;
wire      [9:0] n62;
wire      [9:0] n63;
wire      [9:0] n64;
wire      [9:0] n65;
wire      [9:0] n66;
wire      [9:0] n67;
wire      [9:0] n68;
wire      [9:0] n69;
wire      [9:0] n70;
wire            n71;
wire     [71:0] n72;
wire     [71:0] n73;
wire     [71:0] n74;
wire     [71:0] n75;
wire     [71:0] n76;
wire     [71:0] n77;
wire     [71:0] n78;
wire     [71:0] n79;
wire     [71:0] n80;
wire     [71:0] n81;
wire     [71:0] n82;
wire     [71:0] n83;
wire     [71:0] n84;
wire     [71:0] n85;
wire     [71:0] n86;
wire     [71:0] n87;
wire     [71:0] n88;
wire     [71:0] n89;
wire     [71:0] n90;
wire     [71:0] n91;
wire     [71:0] n92;
wire     [71:0] n93;
wire     [71:0] n94;
wire     [71:0] n95;
wire     [71:0] n96;
wire     [71:0] n97;
wire     [71:0] n98;
wire     [71:0] n99;
wire     [71:0] n100;
wire     [71:0] n101;
wire     [71:0] n102;
wire     [71:0] n103;
wire     [71:0] n104;
wire     [71:0] n105;
wire     [71:0] n106;
wire     [71:0] n107;
wire     [71:0] n108;
wire     [71:0] n109;
wire     [71:0] n110;
wire     [71:0] n111;
wire     [71:0] n112;
wire     [71:0] n113;
wire     [71:0] n114;
wire     [71:0] n115;
wire     [71:0] n116;
wire     [71:0] n117;
wire     [71:0] n118;
wire     [71:0] n119;
wire     [71:0] n120;
wire            n121;
wire      [8:0] n122;
wire      [8:0] n123;
wire      [8:0] n124;
wire      [8:0] n125;
wire      [8:0] n126;
wire      [8:0] n127;
wire      [8:0] n128;
wire      [8:0] n129;
wire            n130;
wire      [9:0] n131;
wire      [9:0] n132;
wire      [9:0] n133;
wire      [9:0] n134;
wire      [9:0] n135;
wire      [9:0] n136;
wire      [9:0] n137;
wire      [9:0] n138;
wire      [9:0] n139;
wire            n140;
wire    [647:0] n141;
wire      [7:0] n142;
wire      [7:0] n143;
wire      [7:0] n144;
wire      [7:0] n145;
wire      [7:0] n146;
wire      [7:0] n147;
wire      [7:0] n148;
wire            n149;
wire            n150;
wire            n151;
wire            n152;
wire            n153;
wire            n154;
wire            n155;
wire            n156;
wire     [18:0] n157;
wire            n158;
wire            n159;
wire            n160;
wire            n161;
wire            n162;
wire            n163;
wire            n164;
wire            n165;
wire     [18:0] n166;
wire            n167;
wire            n168;
wire            n169;
wire            n170;
wire            n171;
wire            n172;
wire            n173;
wire            n174;
wire            n175;
wire            n176;
wire            n177;
wire     [18:0] n178;
wire     [18:0] n179;
wire            n180;
wire            n181;
wire            n182;
wire            n183;
wire            n184;
wire            n185;
wire            n186;
wire            n187;
wire            n188;
wire      [7:0] n189;
wire      [7:0] n190;
wire      [7:0] n191;
wire      [7:0] n192;
wire      [7:0] n193;
wire      [7:0] n194;
wire      [7:0] n195;
wire      [7:0] n196;
wire      [7:0] n197;
wire      [7:0] n198;
wire      [7:0] n199;
wire      [7:0] n200;
wire            n201;
wire            n202;
wire            n203;
wire            n204;
wire            n205;
wire            n206;
wire            n207;
wire            n208;
wire            n209;
wire            n210;
wire            n211;
wire            n212;
wire            n213;
wire            n214;
wire            n215;
wire            n216;
wire      [7:0] n217;
wire            n218;
wire      [7:0] n219;
wire            n220;
wire      [7:0] n221;
wire            n222;
wire      [7:0] n223;
wire            n224;
wire      [7:0] n225;
wire            n226;
wire      [7:0] n227;
wire            n228;
wire      [7:0] n229;
wire            n230;
wire      [7:0] n231;
wire      [7:0] n232;
wire      [7:0] n233;
wire      [7:0] n234;
wire      [7:0] n235;
wire      [7:0] n236;
wire      [7:0] n237;
wire      [7:0] n238;
wire      [7:0] n239;
wire      [7:0] n240;
wire      [7:0] n241;
wire      [7:0] n242;
wire      [7:0] n243;
wire      [7:0] n244;
wire      [7:0] n245;
wire      [7:0] n246;
wire      [7:0] n247;
wire      [7:0] n248;
wire      [7:0] n249;
wire      [7:0] n250;
wire      [7:0] n251;
wire      [7:0] n252;
wire      [7:0] n253;
wire      [7:0] n254;
wire      [7:0] n255;
wire      [7:0] n256;
wire      [7:0] n257;
wire      [7:0] n258;
wire      [7:0] n259;
wire      [7:0] n260;
wire      [7:0] n261;
wire      [7:0] n262;
wire      [7:0] n263;
wire      [7:0] n264;
wire      [7:0] n265;
wire      [7:0] n266;
wire      [7:0] n267;
wire      [7:0] n268;
wire      [7:0] n269;
wire      [7:0] n270;
wire      [7:0] n271;
wire      [7:0] n272;
wire      [7:0] n273;
wire      [7:0] n274;
wire      [7:0] n275;
wire      [7:0] n276;
wire      [7:0] n277;
wire      [7:0] n278;
wire      [7:0] n279;
wire      [7:0] n280;
wire      [7:0] n281;
wire      [7:0] n282;
wire      [7:0] n283;
wire      [7:0] n284;
wire      [7:0] n285;
wire      [7:0] n286;
wire      [7:0] n287;
wire      [7:0] n288;
wire     [15:0] n289;
wire     [23:0] n290;
wire     [31:0] n291;
wire     [39:0] n292;
wire     [47:0] n293;
wire     [55:0] n294;
wire     [63:0] n295;
wire     [71:0] n296;
wire     [71:0] n297;
wire     [71:0] n298;
wire     [71:0] n299;
wire     [71:0] n300;
wire     [71:0] n301;
wire     [71:0] n302;
wire     [71:0] n303;
wire     [71:0] n304;
wire     [71:0] n305;
wire     [71:0] n306;
wire     [71:0] n307;
wire     [71:0] n308;
wire     [71:0] n309;
wire     [71:0] n310;
wire            n311;
wire            n312;
wire            n313;
wire            n314;
wire            n315;
wire            n316;
wire            n317;
wire            n318;
wire            n319;
wire            n320;
wire            n321;
wire            n322;
wire            n323;
wire            n324;
wire            n325;
wire            n326;
wire            n327;
wire            n328;
wire      [7:0] n329;
wire      [7:0] n330;
wire      [7:0] n331;
wire      [7:0] n332;
wire      [7:0] n333;
wire      [7:0] n334;
wire      [7:0] n335;
wire      [7:0] n336;
wire      [7:0] n337;
wire     [15:0] n338;
wire     [23:0] n339;
wire     [31:0] n340;
wire     [39:0] n341;
wire     [47:0] n342;
wire     [55:0] n343;
wire     [63:0] n344;
wire     [71:0] n345;
wire      [7:0] n346;
wire      [7:0] n347;
wire      [7:0] n348;
wire      [7:0] n349;
wire      [7:0] n350;
wire      [7:0] n351;
wire      [7:0] n352;
wire      [7:0] n353;
wire      [7:0] n354;
wire     [15:0] n355;
wire     [23:0] n356;
wire     [31:0] n357;
wire     [39:0] n358;
wire     [47:0] n359;
wire     [55:0] n360;
wire     [63:0] n361;
wire     [71:0] n362;
wire      [7:0] n363;
wire      [7:0] n364;
wire      [7:0] n365;
wire      [7:0] n366;
wire      [7:0] n367;
wire      [7:0] n368;
wire      [7:0] n369;
wire      [7:0] n370;
wire      [7:0] n371;
wire     [15:0] n372;
wire     [23:0] n373;
wire     [31:0] n374;
wire     [39:0] n375;
wire     [47:0] n376;
wire     [55:0] n377;
wire     [63:0] n378;
wire     [71:0] n379;
wire      [7:0] n380;
wire      [7:0] n381;
wire      [7:0] n382;
wire      [7:0] n383;
wire      [7:0] n384;
wire      [7:0] n385;
wire      [7:0] n386;
wire      [7:0] n387;
wire      [7:0] n388;
wire     [15:0] n389;
wire     [23:0] n390;
wire     [31:0] n391;
wire     [39:0] n392;
wire     [47:0] n393;
wire     [55:0] n394;
wire     [63:0] n395;
wire     [71:0] n396;
wire      [7:0] n397;
wire      [7:0] n398;
wire      [7:0] n399;
wire      [7:0] n400;
wire      [7:0] n401;
wire      [7:0] n402;
wire      [7:0] n403;
wire      [7:0] n404;
wire      [7:0] n405;
wire     [15:0] n406;
wire     [23:0] n407;
wire     [31:0] n408;
wire     [39:0] n409;
wire     [47:0] n410;
wire     [55:0] n411;
wire     [63:0] n412;
wire     [71:0] n413;
wire      [7:0] n414;
wire      [7:0] n415;
wire      [7:0] n416;
wire      [7:0] n417;
wire      [7:0] n418;
wire      [7:0] n419;
wire      [7:0] n420;
wire      [7:0] n421;
wire      [7:0] n422;
wire     [15:0] n423;
wire     [23:0] n424;
wire     [31:0] n425;
wire     [39:0] n426;
wire     [47:0] n427;
wire     [55:0] n428;
wire     [63:0] n429;
wire     [71:0] n430;
wire      [7:0] n431;
wire      [7:0] n432;
wire      [7:0] n433;
wire      [7:0] n434;
wire      [7:0] n435;
wire      [7:0] n436;
wire      [7:0] n437;
wire      [7:0] n438;
wire      [7:0] n439;
wire     [15:0] n440;
wire     [23:0] n441;
wire     [31:0] n442;
wire     [39:0] n443;
wire     [47:0] n444;
wire     [55:0] n445;
wire     [63:0] n446;
wire     [71:0] n447;
wire      [7:0] n448;
wire      [7:0] n449;
wire      [7:0] n450;
wire      [7:0] n451;
wire      [7:0] n452;
wire      [7:0] n453;
wire      [7:0] n454;
wire      [7:0] n455;
wire      [7:0] n456;
wire     [15:0] n457;
wire     [23:0] n458;
wire     [31:0] n459;
wire     [39:0] n460;
wire     [47:0] n461;
wire     [55:0] n462;
wire     [63:0] n463;
wire     [71:0] n464;
wire      [7:0] n465;
wire      [7:0] n466;
wire      [7:0] n467;
wire      [7:0] n468;
wire      [7:0] n469;
wire      [7:0] n470;
wire      [7:0] n471;
wire      [7:0] n472;
wire      [7:0] n473;
wire     [15:0] n474;
wire     [23:0] n475;
wire     [31:0] n476;
wire     [39:0] n477;
wire     [47:0] n478;
wire     [55:0] n479;
wire     [63:0] n480;
wire     [71:0] n481;
wire    [143:0] n482;
wire    [215:0] n483;
wire    [287:0] n484;
wire    [359:0] n485;
wire    [431:0] n486;
wire    [503:0] n487;
wire    [575:0] n488;
wire    [647:0] n489;
wire    [647:0] n490;
wire    [647:0] n491;
wire    [647:0] n492;
wire    [647:0] n493;
wire    [647:0] n494;
wire    [647:0] n495;
wire    [647:0] n496;
wire    [647:0] n497;
wire    [647:0] n498;
wire    [647:0] n499;
wire    [647:0] n500;
wire    [647:0] n501;
wire    [647:0] n502;
wire            n503;
wire            n504;
wire            n505;
wire            n506;
wire            n507;
wire            n508;
wire            n509;
wire            n510;
wire            n511;
wire            n512;
wire            n513;
wire            n514;
wire            n515;
wire            n516;
wire            n517;
wire            n518;
wire            n519;
wire            n520;
wire      [8:0] LB2D_proc_0_addr0;
wire      [7:0] LB2D_proc_0_data0;
wire            n521;
wire            n522;
wire            n523;
wire            n524;
wire            n525;
wire            n526;
wire            n527;
wire            n528;
wire            n529;
wire            n530;
wire            n531;
wire            n532;
wire            n533;
wire            n534;
wire            n535;
wire            n536;
wire            n537;
wire            n538;
wire            n539;
wire      [8:0] LB2D_proc_1_addr0;
wire      [7:0] LB2D_proc_1_data0;
wire            n540;
wire            n541;
wire            n542;
wire      [8:0] LB2D_proc_2_addr0;
wire      [7:0] LB2D_proc_2_data0;
wire            n543;
wire            n544;
wire            n545;
wire      [8:0] LB2D_proc_3_addr0;
wire      [7:0] LB2D_proc_3_data0;
wire            n546;
wire            n547;
wire            n548;
wire      [8:0] LB2D_proc_4_addr0;
wire      [7:0] LB2D_proc_4_data0;
wire            n549;
wire            n550;
wire            n551;
wire      [8:0] LB2D_proc_5_addr0;
wire      [7:0] LB2D_proc_5_data0;
wire            n552;
wire            n553;
wire            n554;
wire      [8:0] LB2D_proc_6_addr0;
wire      [7:0] LB2D_proc_6_data0;
wire            n555;
wire            n556;
wire            n557;
wire      [8:0] LB2D_proc_7_addr0;
wire      [7:0] LB2D_proc_7_data0;
wire            n558;
wire            n559;
wire            n560;
wire            n561;
reg      [7:0] LB2D_proc_0[511:0];
reg      [7:0] LB2D_proc_1[511:0];
reg      [7:0] LB2D_proc_2[511:0];
reg      [7:0] LB2D_proc_3[511:0];
reg      [7:0] LB2D_proc_4[511:0];
reg      [7:0] LB2D_proc_5[511:0];
reg      [7:0] LB2D_proc_6[511:0];
reg      [7:0] LB2D_proc_7[511:0];
wire clk;
wire rst;
wire step;
assign n0 =  ( arg_0_TREADY ) == ( 1'd1 )  ;
assign n1 =  ( arg_0_TVALID ) == ( 1'd1 )  ;
assign n2 =  ( n0 ) & ( n1 )  ;
assign n3 =  ( arg_1_TVALID ) == ( 1'd0 )  ;
assign n4 =  ( n2 ) & ( n3 )  ;
assign n5 =  ( arg_1_TREADY ) == ( 1'd1 )  ;
assign n6 =  ( arg_1_TVALID ) == ( 1'd1 )  ;
assign n7 =  ( n5 ) & ( n6 )  ;
assign n8 =  ( arg_0_TREADY ) == ( 1'd0 )  ;
assign n9 =  ( n7 ) & ( n8 )  ;
assign n10 =  ( arg_0_TVALID ) == ( 1'd0 )  ;
assign n11 =  ( gb_exit_it_1 ) == ( 1'd0 )  ;
assign n12 =  ( stencil_stream_empty ) == ( 1'd0 )  ;
assign n13 =  ( n11 ) & ( n12 )  ;
assign n14 =  ( gb_exit_it_1 ) == ( 1'd1 )  ;
assign n15 =  ( gb_exit_it_8 ) == ( 1'd0 )  ;
assign n16 =  ( n14 ) & ( n15 )  ;
assign n17 =  ( n13 ) | ( n16 )  ;
assign n18 =  ( n10 ) & ( n17 )  ;
assign n19 =  ( slice_stream_empty ) == ( 1'd0 )  ;
assign n20 =  ( stencil_stream_full ) == ( 1'd0 )  ;
assign n21 =  ( LB2D_shift_x ) < ( 9'd8 )  ;
assign n22 =  ( n20 ) | ( n21 )  ;
assign n23 =  ( n19 ) & ( n22 )  ;
assign n24 =  ( in_stream_empty ) == ( 1'd0 )  ;
assign n25 =  ( slice_stream_full ) == ( 1'd0 )  ;
assign n26 =  ( LB2D_proc_y ) < ( 10'd8 )  ;
assign n27 =  ( n25 ) | ( n26 )  ;
assign n28 =  ( n24 ) & ( n27 )  ;
assign n29 =  ( arg_1_TREADY ) == ( 1'd0 )  ;
assign n30 =  ( in_stream_full ) == ( 1'd0 )  ;
assign n31 =  ( n29 ) & ( n30 )  ;
assign n32 =  ( LB1D_p_cnt ) != ( 19'd316224 )  ;
assign n33 =  ( n31 ) & ( n32 )  ;
assign n34 =  ( n33 ) ? ( LB1D_buff ) : ( LB1D_buff ) ;
assign n35 =  ( n28 ) ? ( LB1D_buff ) : ( n34 ) ;
assign n36 =  ( n23 ) ? ( LB1D_buff ) : ( n35 ) ;
assign n37 =  ( n18 ) ? ( LB1D_buff ) : ( n36 ) ;
assign n38 =  ( n9 ) ? ( arg_1_TDATA ) : ( n37 ) ;
assign n39 =  ( n4 ) ? ( arg_1_TDATA ) : ( n38 ) ;
assign n40 =  ( LB1D_p_cnt ) + ( 19'd1 )  ;
assign n41 =  ( n33 ) ? ( n40 ) : ( LB1D_p_cnt ) ;
assign n42 =  ( LB2D_proc_w ) < ( 64'd7 )  ;
assign n43 =  ( LB2D_proc_x ) < ( 9'd487 )  ;
assign n44 =  ( LB2D_proc_w ) + ( 64'd1 )  ;
assign n45 =  ( n43 ) ? ( LB2D_proc_w ) : ( n44 ) ;
assign n46 =  ( n42 ) ? ( n45 ) : ( 64'd0 ) ;
assign n47 =  ( n33 ) ? ( LB2D_proc_w ) : ( LB2D_proc_w ) ;
assign n48 =  ( n28 ) ? ( n46 ) : ( n47 ) ;
assign n49 =  ( n23 ) ? ( LB2D_proc_w ) : ( n48 ) ;
assign n50 =  ( n18 ) ? ( LB2D_proc_w ) : ( n49 ) ;
assign n51 =  ( n9 ) ? ( LB2D_proc_w ) : ( n50 ) ;
assign n52 =  ( n4 ) ? ( LB2D_proc_w ) : ( n51 ) ;
assign n53 =  ( LB2D_proc_x ) + ( 9'd1 )  ;
assign n54 =  ( n43 ) ? ( n53 ) : ( 9'd0 ) ;
assign n55 =  ( n33 ) ? ( LB2D_proc_x ) : ( LB2D_proc_x ) ;
assign n56 =  ( n28 ) ? ( n54 ) : ( n55 ) ;
assign n57 =  ( n23 ) ? ( LB2D_proc_x ) : ( n56 ) ;
assign n58 =  ( n18 ) ? ( LB2D_proc_x ) : ( n57 ) ;
assign n59 =  ( n9 ) ? ( LB2D_proc_x ) : ( n58 ) ;
assign n60 =  ( n4 ) ? ( LB2D_proc_x ) : ( n59 ) ;
assign n61 =  ( LB2D_proc_y ) < ( 10'd487 )  ;
assign n62 =  ( LB2D_proc_y ) + ( 10'd1 )  ;
assign n63 =  ( n43 ) ? ( LB2D_proc_y ) : ( n62 ) ;
assign n64 =  ( n61 ) ? ( n63 ) : ( 10'd487 ) ;
assign n65 =  ( n33 ) ? ( LB2D_proc_y ) : ( LB2D_proc_y ) ;
assign n66 =  ( n28 ) ? ( n64 ) : ( n65 ) ;
assign n67 =  ( n23 ) ? ( LB2D_proc_y ) : ( n66 ) ;
assign n68 =  ( n18 ) ? ( LB2D_proc_y ) : ( n67 ) ;
assign n69 =  ( n9 ) ? ( LB2D_proc_y ) : ( n68 ) ;
assign n70 =  ( n4 ) ? ( LB2D_proc_y ) : ( n69 ) ;
assign n71 =  ( slice_stream_full ) == ( 1'd1 )  ;
assign n72 =  ( n71 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n73 =  ( n33 ) ? ( LB2D_shift_0 ) : ( LB2D_shift_0 ) ;
assign n74 =  ( n28 ) ? ( LB2D_shift_0 ) : ( n73 ) ;
assign n75 =  ( n23 ) ? ( n72 ) : ( n74 ) ;
assign n76 =  ( n18 ) ? ( LB2D_shift_0 ) : ( n75 ) ;
assign n77 =  ( n9 ) ? ( LB2D_shift_0 ) : ( n76 ) ;
assign n78 =  ( n4 ) ? ( LB2D_shift_0 ) : ( n77 ) ;
assign n79 =  ( n33 ) ? ( LB2D_shift_1 ) : ( LB2D_shift_1 ) ;
assign n80 =  ( n28 ) ? ( LB2D_shift_1 ) : ( n79 ) ;
assign n81 =  ( n23 ) ? ( LB2D_shift_0 ) : ( n80 ) ;
assign n82 =  ( n18 ) ? ( LB2D_shift_1 ) : ( n81 ) ;
assign n83 =  ( n9 ) ? ( LB2D_shift_1 ) : ( n82 ) ;
assign n84 =  ( n4 ) ? ( LB2D_shift_1 ) : ( n83 ) ;
assign n85 =  ( n33 ) ? ( LB2D_shift_2 ) : ( LB2D_shift_2 ) ;
assign n86 =  ( n28 ) ? ( LB2D_shift_2 ) : ( n85 ) ;
assign n87 =  ( n23 ) ? ( LB2D_shift_1 ) : ( n86 ) ;
assign n88 =  ( n18 ) ? ( LB2D_shift_2 ) : ( n87 ) ;
assign n89 =  ( n9 ) ? ( LB2D_shift_2 ) : ( n88 ) ;
assign n90 =  ( n4 ) ? ( LB2D_shift_2 ) : ( n89 ) ;
assign n91 =  ( n33 ) ? ( LB2D_shift_3 ) : ( LB2D_shift_3 ) ;
assign n92 =  ( n28 ) ? ( LB2D_shift_3 ) : ( n91 ) ;
assign n93 =  ( n23 ) ? ( LB2D_shift_2 ) : ( n92 ) ;
assign n94 =  ( n18 ) ? ( LB2D_shift_3 ) : ( n93 ) ;
assign n95 =  ( n9 ) ? ( LB2D_shift_3 ) : ( n94 ) ;
assign n96 =  ( n4 ) ? ( LB2D_shift_3 ) : ( n95 ) ;
assign n97 =  ( n33 ) ? ( LB2D_shift_4 ) : ( LB2D_shift_4 ) ;
assign n98 =  ( n28 ) ? ( LB2D_shift_4 ) : ( n97 ) ;
assign n99 =  ( n23 ) ? ( LB2D_shift_3 ) : ( n98 ) ;
assign n100 =  ( n18 ) ? ( LB2D_shift_4 ) : ( n99 ) ;
assign n101 =  ( n9 ) ? ( LB2D_shift_4 ) : ( n100 ) ;
assign n102 =  ( n4 ) ? ( LB2D_shift_4 ) : ( n101 ) ;
assign n103 =  ( n33 ) ? ( LB2D_shift_5 ) : ( LB2D_shift_5 ) ;
assign n104 =  ( n28 ) ? ( LB2D_shift_5 ) : ( n103 ) ;
assign n105 =  ( n23 ) ? ( LB2D_shift_4 ) : ( n104 ) ;
assign n106 =  ( n18 ) ? ( LB2D_shift_5 ) : ( n105 ) ;
assign n107 =  ( n9 ) ? ( LB2D_shift_5 ) : ( n106 ) ;
assign n108 =  ( n4 ) ? ( LB2D_shift_5 ) : ( n107 ) ;
assign n109 =  ( n33 ) ? ( LB2D_shift_6 ) : ( LB2D_shift_6 ) ;
assign n110 =  ( n28 ) ? ( LB2D_shift_6 ) : ( n109 ) ;
assign n111 =  ( n23 ) ? ( LB2D_shift_5 ) : ( n110 ) ;
assign n112 =  ( n18 ) ? ( LB2D_shift_6 ) : ( n111 ) ;
assign n113 =  ( n9 ) ? ( LB2D_shift_6 ) : ( n112 ) ;
assign n114 =  ( n4 ) ? ( LB2D_shift_6 ) : ( n113 ) ;
assign n115 =  ( n33 ) ? ( LB2D_shift_7 ) : ( LB2D_shift_7 ) ;
assign n116 =  ( n28 ) ? ( LB2D_shift_7 ) : ( n115 ) ;
assign n117 =  ( n23 ) ? ( LB2D_shift_6 ) : ( n116 ) ;
assign n118 =  ( n18 ) ? ( LB2D_shift_7 ) : ( n117 ) ;
assign n119 =  ( n9 ) ? ( LB2D_shift_7 ) : ( n118 ) ;
assign n120 =  ( n4 ) ? ( LB2D_shift_7 ) : ( n119 ) ;
assign n121 =  ( LB2D_shift_x ) < ( 9'd487 )  ;
assign n122 =  ( LB2D_shift_x ) + ( 9'd1 )  ;
assign n123 =  ( n121 ) ? ( n122 ) : ( 9'd0 ) ;
assign n124 =  ( n33 ) ? ( LB2D_shift_x ) : ( LB2D_shift_x ) ;
assign n125 =  ( n28 ) ? ( LB2D_shift_x ) : ( n124 ) ;
assign n126 =  ( n23 ) ? ( n123 ) : ( n125 ) ;
assign n127 =  ( n18 ) ? ( LB2D_shift_x ) : ( n126 ) ;
assign n128 =  ( n9 ) ? ( LB2D_shift_x ) : ( n127 ) ;
assign n129 =  ( n4 ) ? ( LB2D_shift_x ) : ( n128 ) ;
assign n130 =  ( LB2D_shift_y ) < ( 10'd479 )  ;
assign n131 =  ( LB2D_shift_y ) + ( 10'd1 )  ;
assign n132 =  ( n121 ) ? ( LB2D_shift_y ) : ( n131 ) ;
assign n133 =  ( n130 ) ? ( n132 ) : ( 10'd479 ) ;
assign n134 =  ( n33 ) ? ( LB2D_shift_y ) : ( LB2D_shift_y ) ;
assign n135 =  ( n28 ) ? ( LB2D_shift_y ) : ( n134 ) ;
assign n136 =  ( n23 ) ? ( n133 ) : ( n135 ) ;
assign n137 =  ( n18 ) ? ( LB2D_shift_y ) : ( n136 ) ;
assign n138 =  ( n9 ) ? ( LB2D_shift_y ) : ( n137 ) ;
assign n139 =  ( n4 ) ? ( LB2D_shift_y ) : ( n138 ) ;
assign n140 =  ( stencil_stream_full ) == ( 1'd1 )  ;
assign n141 =  ( n140 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_0 ) ;
assign n142 = gb_fun(n141) ;
assign n143 =  ( n33 ) ? ( arg_0_TDATA ) : ( arg_0_TDATA ) ;
assign n144 =  ( n28 ) ? ( arg_0_TDATA ) : ( n143 ) ;
assign n145 =  ( n23 ) ? ( arg_0_TDATA ) : ( n144 ) ;
assign n146 =  ( n18 ) ? ( n142 ) : ( n145 ) ;
assign n147 =  ( n9 ) ? ( arg_0_TDATA ) : ( n146 ) ;
assign n148 =  ( n4 ) ? ( arg_0_TDATA ) : ( n147 ) ;
assign n149 =  ( gb_pp_it_8 ) == ( 1'd1 )  ;
assign n150 =  ( n149 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n151 =  ( n33 ) ? ( arg_0_TVALID ) : ( arg_0_TVALID ) ;
assign n152 =  ( n28 ) ? ( arg_0_TVALID ) : ( n151 ) ;
assign n153 =  ( n23 ) ? ( arg_0_TVALID ) : ( n152 ) ;
assign n154 =  ( n18 ) ? ( n150 ) : ( n153 ) ;
assign n155 =  ( n9 ) ? ( arg_0_TVALID ) : ( n154 ) ;
assign n156 =  ( n4 ) ? ( 1'd0 ) : ( n155 ) ;
assign n157 =  ( 19'd316224 ) - ( 19'd1 )  ;
assign n158 =  ( LB1D_p_cnt ) == ( n157 )  ;
assign n159 =  ( n158 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n160 =  ( n33 ) ? ( n159 ) : ( arg_1_TREADY ) ;
assign n161 =  ( n28 ) ? ( arg_1_TREADY ) : ( n160 ) ;
assign n162 =  ( n23 ) ? ( arg_1_TREADY ) : ( n161 ) ;
assign n163 =  ( n18 ) ? ( arg_1_TREADY ) : ( n162 ) ;
assign n164 =  ( n9 ) ? ( 1'd0 ) : ( n163 ) ;
assign n165 =  ( n4 ) ? ( 1'd0 ) : ( n164 ) ;
assign n166 =  ( gb_p_cnt ) + ( 19'd1 )  ;
assign n167 =  ( n166 ) == ( 19'd307200 )  ;
assign n168 =  ( n167 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n169 =  ( n18 ) ? ( n168 ) : ( gb_exit_it_1 ) ;
assign n170 =  ( n18 ) ? ( gb_exit_it_1 ) : ( gb_exit_it_2 ) ;
assign n171 =  ( n18 ) ? ( gb_exit_it_2 ) : ( gb_exit_it_3 ) ;
assign n172 =  ( n18 ) ? ( gb_exit_it_3 ) : ( gb_exit_it_4 ) ;
assign n173 =  ( n18 ) ? ( gb_exit_it_4 ) : ( gb_exit_it_5 ) ;
assign n174 =  ( n18 ) ? ( gb_exit_it_5 ) : ( gb_exit_it_6 ) ;
assign n175 =  ( n18 ) ? ( gb_exit_it_6 ) : ( gb_exit_it_7 ) ;
assign n176 =  ( n18 ) ? ( gb_exit_it_7 ) : ( gb_exit_it_8 ) ;
assign n177 =  ( gb_p_cnt ) < ( 19'd307200 )  ;
assign n178 =  ( n177 ) ? ( n166 ) : ( 19'd307200 ) ;
assign n179 =  ( n18 ) ? ( n178 ) : ( gb_p_cnt ) ;
assign n180 =  ( n18 ) ? ( 1'd1 ) : ( gb_pp_it_1 ) ;
assign n181 =  ( n18 ) ? ( gb_pp_it_1 ) : ( gb_pp_it_2 ) ;
assign n182 =  ( n18 ) ? ( gb_pp_it_2 ) : ( gb_pp_it_3 ) ;
assign n183 =  ( n18 ) ? ( gb_pp_it_3 ) : ( gb_pp_it_4 ) ;
assign n184 =  ( n18 ) ? ( gb_pp_it_4 ) : ( gb_pp_it_5 ) ;
assign n185 =  ( n18 ) ? ( gb_pp_it_5 ) : ( gb_pp_it_6 ) ;
assign n186 =  ( n18 ) ? ( gb_pp_it_6 ) : ( gb_pp_it_7 ) ;
assign n187 =  ( n18 ) ? ( gb_pp_it_7 ) : ( gb_pp_it_8 ) ;
assign n188 =  ( n18 ) ? ( gb_pp_it_8 ) : ( gb_pp_it_9 ) ;
assign n189 =  ( n33 ) ? ( LB1D_buff ) : ( in_stream_buff_0 ) ;
assign n190 =  ( n28 ) ? ( in_stream_buff_0 ) : ( n189 ) ;
assign n191 =  ( n23 ) ? ( in_stream_buff_0 ) : ( n190 ) ;
assign n192 =  ( n18 ) ? ( in_stream_buff_0 ) : ( n191 ) ;
assign n193 =  ( n9 ) ? ( in_stream_buff_0 ) : ( n192 ) ;
assign n194 =  ( n4 ) ? ( in_stream_buff_0 ) : ( n193 ) ;
assign n195 =  ( n33 ) ? ( in_stream_buff_0 ) : ( in_stream_buff_1 ) ;
assign n196 =  ( n28 ) ? ( in_stream_buff_1 ) : ( n195 ) ;
assign n197 =  ( n23 ) ? ( in_stream_buff_1 ) : ( n196 ) ;
assign n198 =  ( n18 ) ? ( in_stream_buff_1 ) : ( n197 ) ;
assign n199 =  ( n9 ) ? ( in_stream_buff_1 ) : ( n198 ) ;
assign n200 =  ( n4 ) ? ( in_stream_buff_1 ) : ( n199 ) ;
assign n201 =  ( in_stream_full ) == ( 1'd1 )  ;
assign n202 =  ( n201 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n203 =  ( n33 ) ? ( 1'd0 ) : ( in_stream_empty ) ;
assign n204 =  ( n28 ) ? ( n202 ) : ( n203 ) ;
assign n205 =  ( n23 ) ? ( in_stream_empty ) : ( n204 ) ;
assign n206 =  ( n18 ) ? ( in_stream_empty ) : ( n205 ) ;
assign n207 =  ( n9 ) ? ( in_stream_empty ) : ( n206 ) ;
assign n208 =  ( n4 ) ? ( in_stream_empty ) : ( n207 ) ;
assign n209 =  ( in_stream_empty ) == ( 1'd1 )  ;
assign n210 =  ( n209 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n211 =  ( n33 ) ? ( n210 ) : ( in_stream_full ) ;
assign n212 =  ( n28 ) ? ( 1'd0 ) : ( n211 ) ;
assign n213 =  ( n23 ) ? ( in_stream_full ) : ( n212 ) ;
assign n214 =  ( n18 ) ? ( in_stream_full ) : ( n213 ) ;
assign n215 =  ( n9 ) ? ( in_stream_full ) : ( n214 ) ;
assign n216 =  ( n4 ) ? ( in_stream_full ) : ( n215 ) ;
assign n217 =  ( n201 ) ? ( in_stream_buff_1 ) : ( in_stream_buff_0 ) ;
assign n218 =  ( LB2D_proc_w ) == ( 64'd0 )  ;
assign n219 =  (  LB2D_proc_7 [ LB2D_proc_x ] )  ;
assign n220 =  ( LB2D_proc_w ) == ( 64'd1 )  ;
assign n221 =  (  LB2D_proc_0 [ LB2D_proc_x ] )  ;
assign n222 =  ( LB2D_proc_w ) == ( 64'd2 )  ;
assign n223 =  (  LB2D_proc_1 [ LB2D_proc_x ] )  ;
assign n224 =  ( LB2D_proc_w ) == ( 64'd3 )  ;
assign n225 =  (  LB2D_proc_2 [ LB2D_proc_x ] )  ;
assign n226 =  ( LB2D_proc_w ) == ( 64'd4 )  ;
assign n227 =  (  LB2D_proc_3 [ LB2D_proc_x ] )  ;
assign n228 =  ( LB2D_proc_w ) == ( 64'd5 )  ;
assign n229 =  (  LB2D_proc_4 [ LB2D_proc_x ] )  ;
assign n230 =  ( LB2D_proc_w ) == ( 64'd6 )  ;
assign n231 =  (  LB2D_proc_5 [ LB2D_proc_x ] )  ;
assign n232 =  (  LB2D_proc_6 [ LB2D_proc_x ] )  ;
assign n233 =  ( n230 ) ? ( n231 ) : ( n232 ) ;
assign n234 =  ( n228 ) ? ( n229 ) : ( n233 ) ;
assign n235 =  ( n226 ) ? ( n227 ) : ( n234 ) ;
assign n236 =  ( n224 ) ? ( n225 ) : ( n235 ) ;
assign n237 =  ( n222 ) ? ( n223 ) : ( n236 ) ;
assign n238 =  ( n220 ) ? ( n221 ) : ( n237 ) ;
assign n239 =  ( n218 ) ? ( n219 ) : ( n238 ) ;
assign n240 =  ( n230 ) ? ( n229 ) : ( n231 ) ;
assign n241 =  ( n228 ) ? ( n227 ) : ( n240 ) ;
assign n242 =  ( n226 ) ? ( n225 ) : ( n241 ) ;
assign n243 =  ( n224 ) ? ( n223 ) : ( n242 ) ;
assign n244 =  ( n222 ) ? ( n221 ) : ( n243 ) ;
assign n245 =  ( n220 ) ? ( n219 ) : ( n244 ) ;
assign n246 =  ( n218 ) ? ( n232 ) : ( n245 ) ;
assign n247 =  ( n230 ) ? ( n227 ) : ( n229 ) ;
assign n248 =  ( n228 ) ? ( n225 ) : ( n247 ) ;
assign n249 =  ( n226 ) ? ( n223 ) : ( n248 ) ;
assign n250 =  ( n224 ) ? ( n221 ) : ( n249 ) ;
assign n251 =  ( n222 ) ? ( n219 ) : ( n250 ) ;
assign n252 =  ( n220 ) ? ( n232 ) : ( n251 ) ;
assign n253 =  ( n218 ) ? ( n231 ) : ( n252 ) ;
assign n254 =  ( n230 ) ? ( n225 ) : ( n227 ) ;
assign n255 =  ( n228 ) ? ( n223 ) : ( n254 ) ;
assign n256 =  ( n226 ) ? ( n221 ) : ( n255 ) ;
assign n257 =  ( n224 ) ? ( n219 ) : ( n256 ) ;
assign n258 =  ( n222 ) ? ( n232 ) : ( n257 ) ;
assign n259 =  ( n220 ) ? ( n231 ) : ( n258 ) ;
assign n260 =  ( n218 ) ? ( n229 ) : ( n259 ) ;
assign n261 =  ( n230 ) ? ( n223 ) : ( n225 ) ;
assign n262 =  ( n228 ) ? ( n221 ) : ( n261 ) ;
assign n263 =  ( n226 ) ? ( n219 ) : ( n262 ) ;
assign n264 =  ( n224 ) ? ( n232 ) : ( n263 ) ;
assign n265 =  ( n222 ) ? ( n231 ) : ( n264 ) ;
assign n266 =  ( n220 ) ? ( n229 ) : ( n265 ) ;
assign n267 =  ( n218 ) ? ( n227 ) : ( n266 ) ;
assign n268 =  ( n230 ) ? ( n221 ) : ( n223 ) ;
assign n269 =  ( n228 ) ? ( n219 ) : ( n268 ) ;
assign n270 =  ( n226 ) ? ( n232 ) : ( n269 ) ;
assign n271 =  ( n224 ) ? ( n231 ) : ( n270 ) ;
assign n272 =  ( n222 ) ? ( n229 ) : ( n271 ) ;
assign n273 =  ( n220 ) ? ( n227 ) : ( n272 ) ;
assign n274 =  ( n218 ) ? ( n225 ) : ( n273 ) ;
assign n275 =  ( n230 ) ? ( n219 ) : ( n221 ) ;
assign n276 =  ( n228 ) ? ( n232 ) : ( n275 ) ;
assign n277 =  ( n226 ) ? ( n231 ) : ( n276 ) ;
assign n278 =  ( n224 ) ? ( n229 ) : ( n277 ) ;
assign n279 =  ( n222 ) ? ( n227 ) : ( n278 ) ;
assign n280 =  ( n220 ) ? ( n225 ) : ( n279 ) ;
assign n281 =  ( n218 ) ? ( n223 ) : ( n280 ) ;
assign n282 =  ( n230 ) ? ( n232 ) : ( n219 ) ;
assign n283 =  ( n228 ) ? ( n231 ) : ( n282 ) ;
assign n284 =  ( n226 ) ? ( n229 ) : ( n283 ) ;
assign n285 =  ( n224 ) ? ( n227 ) : ( n284 ) ;
assign n286 =  ( n222 ) ? ( n225 ) : ( n285 ) ;
assign n287 =  ( n220 ) ? ( n223 ) : ( n286 ) ;
assign n288 =  ( n218 ) ? ( n221 ) : ( n287 ) ;
assign n289 =  { ( n281 ) , ( n288 ) }  ;
assign n290 =  { ( n274 ) , ( n289 ) }  ;
assign n291 =  { ( n267 ) , ( n290 ) }  ;
assign n292 =  { ( n260 ) , ( n291 ) }  ;
assign n293 =  { ( n253 ) , ( n292 ) }  ;
assign n294 =  { ( n246 ) , ( n293 ) }  ;
assign n295 =  { ( n239 ) , ( n294 ) }  ;
assign n296 =  { ( n217 ) , ( n295 ) }  ;
assign n297 =  ( n26 ) ? ( slice_stream_buff_0 ) : ( n296 ) ;
assign n298 =  ( n33 ) ? ( slice_stream_buff_0 ) : ( slice_stream_buff_0 ) ;
assign n299 =  ( n28 ) ? ( n297 ) : ( n298 ) ;
assign n300 =  ( n23 ) ? ( slice_stream_buff_0 ) : ( n299 ) ;
assign n301 =  ( n18 ) ? ( slice_stream_buff_0 ) : ( n300 ) ;
assign n302 =  ( n9 ) ? ( slice_stream_buff_0 ) : ( n301 ) ;
assign n303 =  ( n4 ) ? ( slice_stream_buff_0 ) : ( n302 ) ;
assign n304 =  ( n26 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n305 =  ( n33 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_1 ) ;
assign n306 =  ( n28 ) ? ( n304 ) : ( n305 ) ;
assign n307 =  ( n23 ) ? ( slice_stream_buff_1 ) : ( n306 ) ;
assign n308 =  ( n18 ) ? ( slice_stream_buff_1 ) : ( n307 ) ;
assign n309 =  ( n9 ) ? ( slice_stream_buff_1 ) : ( n308 ) ;
assign n310 =  ( n4 ) ? ( slice_stream_buff_1 ) : ( n309 ) ;
assign n311 =  ( n71 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n312 =  ( n26 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n313 =  ( n33 ) ? ( slice_stream_empty ) : ( slice_stream_empty ) ;
assign n314 =  ( n28 ) ? ( n312 ) : ( n313 ) ;
assign n315 =  ( n23 ) ? ( n311 ) : ( n314 ) ;
assign n316 =  ( n18 ) ? ( slice_stream_empty ) : ( n315 ) ;
assign n317 =  ( n9 ) ? ( slice_stream_empty ) : ( n316 ) ;
assign n318 =  ( n4 ) ? ( slice_stream_empty ) : ( n317 ) ;
assign n319 =  ( slice_stream_empty ) == ( 1'd1 )  ;
assign n320 =  ( n319 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n321 =  ( n26 ) ? ( 1'd0 ) : ( n320 ) ;
assign n322 =  ( n33 ) ? ( slice_stream_full ) : ( slice_stream_full ) ;
assign n323 =  ( n28 ) ? ( n321 ) : ( n322 ) ;
assign n324 =  ( n23 ) ? ( 1'd0 ) : ( n323 ) ;
assign n325 =  ( n18 ) ? ( slice_stream_full ) : ( n324 ) ;
assign n326 =  ( n9 ) ? ( slice_stream_full ) : ( n325 ) ;
assign n327 =  ( n4 ) ? ( slice_stream_full ) : ( n326 ) ;
assign n328 =  ( LB2D_shift_x ) >= ( 9'd8 )  ;
assign n329 = n72[71:64] ;
assign n330 = LB2D_shift_0[71:64] ;
assign n331 = LB2D_shift_1[71:64] ;
assign n332 = LB2D_shift_2[71:64] ;
assign n333 = LB2D_shift_3[71:64] ;
assign n334 = LB2D_shift_4[71:64] ;
assign n335 = LB2D_shift_5[71:64] ;
assign n336 = LB2D_shift_6[71:64] ;
assign n337 = LB2D_shift_7[71:64] ;
assign n338 =  { ( n336 ) , ( n337 ) }  ;
assign n339 =  { ( n335 ) , ( n338 ) }  ;
assign n340 =  { ( n334 ) , ( n339 ) }  ;
assign n341 =  { ( n333 ) , ( n340 ) }  ;
assign n342 =  { ( n332 ) , ( n341 ) }  ;
assign n343 =  { ( n331 ) , ( n342 ) }  ;
assign n344 =  { ( n330 ) , ( n343 ) }  ;
assign n345 =  { ( n329 ) , ( n344 ) }  ;
assign n346 = n72[63:56] ;
assign n347 = LB2D_shift_0[63:56] ;
assign n348 = LB2D_shift_1[63:56] ;
assign n349 = LB2D_shift_2[63:56] ;
assign n350 = LB2D_shift_3[63:56] ;
assign n351 = LB2D_shift_4[63:56] ;
assign n352 = LB2D_shift_5[63:56] ;
assign n353 = LB2D_shift_6[63:56] ;
assign n354 = LB2D_shift_7[63:56] ;
assign n355 =  { ( n353 ) , ( n354 ) }  ;
assign n356 =  { ( n352 ) , ( n355 ) }  ;
assign n357 =  { ( n351 ) , ( n356 ) }  ;
assign n358 =  { ( n350 ) , ( n357 ) }  ;
assign n359 =  { ( n349 ) , ( n358 ) }  ;
assign n360 =  { ( n348 ) , ( n359 ) }  ;
assign n361 =  { ( n347 ) , ( n360 ) }  ;
assign n362 =  { ( n346 ) , ( n361 ) }  ;
assign n363 = n72[55:48] ;
assign n364 = LB2D_shift_0[55:48] ;
assign n365 = LB2D_shift_1[55:48] ;
assign n366 = LB2D_shift_2[55:48] ;
assign n367 = LB2D_shift_3[55:48] ;
assign n368 = LB2D_shift_4[55:48] ;
assign n369 = LB2D_shift_5[55:48] ;
assign n370 = LB2D_shift_6[55:48] ;
assign n371 = LB2D_shift_7[55:48] ;
assign n372 =  { ( n370 ) , ( n371 ) }  ;
assign n373 =  { ( n369 ) , ( n372 ) }  ;
assign n374 =  { ( n368 ) , ( n373 ) }  ;
assign n375 =  { ( n367 ) , ( n374 ) }  ;
assign n376 =  { ( n366 ) , ( n375 ) }  ;
assign n377 =  { ( n365 ) , ( n376 ) }  ;
assign n378 =  { ( n364 ) , ( n377 ) }  ;
assign n379 =  { ( n363 ) , ( n378 ) }  ;
assign n380 = n72[47:40] ;
assign n381 = LB2D_shift_0[47:40] ;
assign n382 = LB2D_shift_1[47:40] ;
assign n383 = LB2D_shift_2[47:40] ;
assign n384 = LB2D_shift_3[47:40] ;
assign n385 = LB2D_shift_4[47:40] ;
assign n386 = LB2D_shift_5[47:40] ;
assign n387 = LB2D_shift_6[47:40] ;
assign n388 = LB2D_shift_7[47:40] ;
assign n389 =  { ( n387 ) , ( n388 ) }  ;
assign n390 =  { ( n386 ) , ( n389 ) }  ;
assign n391 =  { ( n385 ) , ( n390 ) }  ;
assign n392 =  { ( n384 ) , ( n391 ) }  ;
assign n393 =  { ( n383 ) , ( n392 ) }  ;
assign n394 =  { ( n382 ) , ( n393 ) }  ;
assign n395 =  { ( n381 ) , ( n394 ) }  ;
assign n396 =  { ( n380 ) , ( n395 ) }  ;
assign n397 = n72[39:32] ;
assign n398 = LB2D_shift_0[39:32] ;
assign n399 = LB2D_shift_1[39:32] ;
assign n400 = LB2D_shift_2[39:32] ;
assign n401 = LB2D_shift_3[39:32] ;
assign n402 = LB2D_shift_4[39:32] ;
assign n403 = LB2D_shift_5[39:32] ;
assign n404 = LB2D_shift_6[39:32] ;
assign n405 = LB2D_shift_7[39:32] ;
assign n406 =  { ( n404 ) , ( n405 ) }  ;
assign n407 =  { ( n403 ) , ( n406 ) }  ;
assign n408 =  { ( n402 ) , ( n407 ) }  ;
assign n409 =  { ( n401 ) , ( n408 ) }  ;
assign n410 =  { ( n400 ) , ( n409 ) }  ;
assign n411 =  { ( n399 ) , ( n410 ) }  ;
assign n412 =  { ( n398 ) , ( n411 ) }  ;
assign n413 =  { ( n397 ) , ( n412 ) }  ;
assign n414 = n72[31:24] ;
assign n415 = LB2D_shift_0[31:24] ;
assign n416 = LB2D_shift_1[31:24] ;
assign n417 = LB2D_shift_2[31:24] ;
assign n418 = LB2D_shift_3[31:24] ;
assign n419 = LB2D_shift_4[31:24] ;
assign n420 = LB2D_shift_5[31:24] ;
assign n421 = LB2D_shift_6[31:24] ;
assign n422 = LB2D_shift_7[31:24] ;
assign n423 =  { ( n421 ) , ( n422 ) }  ;
assign n424 =  { ( n420 ) , ( n423 ) }  ;
assign n425 =  { ( n419 ) , ( n424 ) }  ;
assign n426 =  { ( n418 ) , ( n425 ) }  ;
assign n427 =  { ( n417 ) , ( n426 ) }  ;
assign n428 =  { ( n416 ) , ( n427 ) }  ;
assign n429 =  { ( n415 ) , ( n428 ) }  ;
assign n430 =  { ( n414 ) , ( n429 ) }  ;
assign n431 = n72[23:16] ;
assign n432 = LB2D_shift_0[23:16] ;
assign n433 = LB2D_shift_1[23:16] ;
assign n434 = LB2D_shift_2[23:16] ;
assign n435 = LB2D_shift_3[23:16] ;
assign n436 = LB2D_shift_4[23:16] ;
assign n437 = LB2D_shift_5[23:16] ;
assign n438 = LB2D_shift_6[23:16] ;
assign n439 = LB2D_shift_7[23:16] ;
assign n440 =  { ( n438 ) , ( n439 ) }  ;
assign n441 =  { ( n437 ) , ( n440 ) }  ;
assign n442 =  { ( n436 ) , ( n441 ) }  ;
assign n443 =  { ( n435 ) , ( n442 ) }  ;
assign n444 =  { ( n434 ) , ( n443 ) }  ;
assign n445 =  { ( n433 ) , ( n444 ) }  ;
assign n446 =  { ( n432 ) , ( n445 ) }  ;
assign n447 =  { ( n431 ) , ( n446 ) }  ;
assign n448 = n72[15:8] ;
assign n449 = LB2D_shift_0[15:8] ;
assign n450 = LB2D_shift_1[15:8] ;
assign n451 = LB2D_shift_2[15:8] ;
assign n452 = LB2D_shift_3[15:8] ;
assign n453 = LB2D_shift_4[15:8] ;
assign n454 = LB2D_shift_5[15:8] ;
assign n455 = LB2D_shift_6[15:8] ;
assign n456 = LB2D_shift_7[15:8] ;
assign n457 =  { ( n455 ) , ( n456 ) }  ;
assign n458 =  { ( n454 ) , ( n457 ) }  ;
assign n459 =  { ( n453 ) , ( n458 ) }  ;
assign n460 =  { ( n452 ) , ( n459 ) }  ;
assign n461 =  { ( n451 ) , ( n460 ) }  ;
assign n462 =  { ( n450 ) , ( n461 ) }  ;
assign n463 =  { ( n449 ) , ( n462 ) }  ;
assign n464 =  { ( n448 ) , ( n463 ) }  ;
assign n465 = n72[7:0] ;
assign n466 = LB2D_shift_0[7:0] ;
assign n467 = LB2D_shift_1[7:0] ;
assign n468 = LB2D_shift_2[7:0] ;
assign n469 = LB2D_shift_3[7:0] ;
assign n470 = LB2D_shift_4[7:0] ;
assign n471 = LB2D_shift_5[7:0] ;
assign n472 = LB2D_shift_6[7:0] ;
assign n473 = LB2D_shift_7[7:0] ;
assign n474 =  { ( n472 ) , ( n473 ) }  ;
assign n475 =  { ( n471 ) , ( n474 ) }  ;
assign n476 =  { ( n470 ) , ( n475 ) }  ;
assign n477 =  { ( n469 ) , ( n476 ) }  ;
assign n478 =  { ( n468 ) , ( n477 ) }  ;
assign n479 =  { ( n467 ) , ( n478 ) }  ;
assign n480 =  { ( n466 ) , ( n479 ) }  ;
assign n481 =  { ( n465 ) , ( n480 ) }  ;
assign n482 =  { ( n464 ) , ( n481 ) }  ;
assign n483 =  { ( n447 ) , ( n482 ) }  ;
assign n484 =  { ( n430 ) , ( n483 ) }  ;
assign n485 =  { ( n413 ) , ( n484 ) }  ;
assign n486 =  { ( n396 ) , ( n485 ) }  ;
assign n487 =  { ( n379 ) , ( n486 ) }  ;
assign n488 =  { ( n362 ) , ( n487 ) }  ;
assign n489 =  { ( n345 ) , ( n488 ) }  ;
assign n490 =  ( n328 ) ? ( n489 ) : ( stencil_stream_buff_0 ) ;
assign n491 =  ( n33 ) ? ( stencil_stream_buff_0 ) : ( stencil_stream_buff_0 ) ;
assign n492 =  ( n28 ) ? ( stencil_stream_buff_0 ) : ( n491 ) ;
assign n493 =  ( n23 ) ? ( n490 ) : ( n492 ) ;
assign n494 =  ( n18 ) ? ( stencil_stream_buff_0 ) : ( n493 ) ;
assign n495 =  ( n9 ) ? ( stencil_stream_buff_0 ) : ( n494 ) ;
assign n496 =  ( n4 ) ? ( stencil_stream_buff_0 ) : ( n495 ) ;
assign n497 =  ( n33 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_1 ) ;
assign n498 =  ( n28 ) ? ( stencil_stream_buff_1 ) : ( n497 ) ;
assign n499 =  ( n23 ) ? ( stencil_stream_buff_0 ) : ( n498 ) ;
assign n500 =  ( n18 ) ? ( stencil_stream_buff_1 ) : ( n499 ) ;
assign n501 =  ( n9 ) ? ( stencil_stream_buff_1 ) : ( n500 ) ;
assign n502 =  ( n4 ) ? ( stencil_stream_buff_1 ) : ( n501 ) ;
assign n503 =  ( n140 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n504 =  ( n21 ) ? ( stencil_stream_empty ) : ( 1'd0 ) ;
assign n505 =  ( n33 ) ? ( stencil_stream_empty ) : ( stencil_stream_empty ) ;
assign n506 =  ( n28 ) ? ( stencil_stream_empty ) : ( n505 ) ;
assign n507 =  ( n23 ) ? ( n504 ) : ( n506 ) ;
assign n508 =  ( n18 ) ? ( n503 ) : ( n507 ) ;
assign n509 =  ( n9 ) ? ( stencil_stream_empty ) : ( n508 ) ;
assign n510 =  ( n4 ) ? ( stencil_stream_empty ) : ( n509 ) ;
assign n511 =  ( n14 ) ? ( 1'd0 ) : ( 1'd0 ) ;
assign n512 =  ( stencil_stream_empty ) == ( 1'd1 )  ;
assign n513 =  ( n512 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n514 =  ( n21 ) ? ( stencil_stream_full ) : ( n513 ) ;
assign n515 =  ( n33 ) ? ( stencil_stream_full ) : ( stencil_stream_full ) ;
assign n516 =  ( n28 ) ? ( stencil_stream_full ) : ( n515 ) ;
assign n517 =  ( n23 ) ? ( n514 ) : ( n516 ) ;
assign n518 =  ( n18 ) ? ( n511 ) : ( n517 ) ;
assign n519 =  ( n9 ) ? ( stencil_stream_full ) : ( n518 ) ;
assign n520 =  ( n4 ) ? ( stencil_stream_full ) : ( n519 ) ;
assign n521 = ~ ( n4 ) ;
assign n522 = ~ ( n9 ) ;
assign n523 =  ( n521 ) & ( n522 )  ;
assign n524 = ~ ( n18 ) ;
assign n525 =  ( n523 ) & ( n524 )  ;
assign n526 = ~ ( n23 ) ;
assign n527 =  ( n525 ) & ( n526 )  ;
assign n528 = ~ ( n28 ) ;
assign n529 =  ( n527 ) & ( n528 )  ;
assign n530 = ~ ( n33 ) ;
assign n531 =  ( n529 ) & ( n530 )  ;
assign n532 =  ( n529 ) & ( n33 )  ;
assign n533 =  ( n527 ) & ( n28 )  ;
assign n534 = ~ ( n218 ) ;
assign n535 =  ( n533 ) & ( n534 )  ;
assign n536 =  ( n533 ) & ( n218 )  ;
assign n537 =  ( n525 ) & ( n23 )  ;
assign n538 =  ( n523 ) & ( n18 )  ;
assign n539 =  ( n521 ) & ( n9 )  ;
assign LB2D_proc_0_addr0 = n536 ? (LB2D_proc_x) : (0);
assign LB2D_proc_0_data0 = n536 ? (n217) : (LB2D_proc_0[0]);
assign n540 = ~ ( n220 ) ;
assign n541 =  ( n533 ) & ( n540 )  ;
assign n542 =  ( n533 ) & ( n220 )  ;
assign LB2D_proc_1_addr0 = n542 ? (LB2D_proc_x) : (0);
assign LB2D_proc_1_data0 = n542 ? (n217) : (LB2D_proc_1[0]);
assign n543 = ~ ( n222 ) ;
assign n544 =  ( n533 ) & ( n543 )  ;
assign n545 =  ( n533 ) & ( n222 )  ;
assign LB2D_proc_2_addr0 = n545 ? (LB2D_proc_x) : (0);
assign LB2D_proc_2_data0 = n545 ? (n217) : (LB2D_proc_2[0]);
assign n546 = ~ ( n224 ) ;
assign n547 =  ( n533 ) & ( n546 )  ;
assign n548 =  ( n533 ) & ( n224 )  ;
assign LB2D_proc_3_addr0 = n548 ? (LB2D_proc_x) : (0);
assign LB2D_proc_3_data0 = n548 ? (n217) : (LB2D_proc_3[0]);
assign n549 = ~ ( n226 ) ;
assign n550 =  ( n533 ) & ( n549 )  ;
assign n551 =  ( n533 ) & ( n226 )  ;
assign LB2D_proc_4_addr0 = n551 ? (LB2D_proc_x) : (0);
assign LB2D_proc_4_data0 = n551 ? (n217) : (LB2D_proc_4[0]);
assign n552 = ~ ( n228 ) ;
assign n553 =  ( n533 ) & ( n552 )  ;
assign n554 =  ( n533 ) & ( n228 )  ;
assign LB2D_proc_5_addr0 = n554 ? (LB2D_proc_x) : (0);
assign LB2D_proc_5_data0 = n554 ? (n217) : (LB2D_proc_5[0]);
assign n555 = ~ ( n230 ) ;
assign n556 =  ( n533 ) & ( n555 )  ;
assign n557 =  ( n533 ) & ( n230 )  ;
assign LB2D_proc_6_addr0 = n557 ? (LB2D_proc_x) : (0);
assign LB2D_proc_6_data0 = n557 ? (n217) : (LB2D_proc_6[0]);
assign n558 =  ( LB2D_proc_w ) == ( 64'd7 )  ;
assign n559 = ~ ( n558 ) ;
assign n560 =  ( n533 ) & ( n559 )  ;
assign n561 =  ( n533 ) & ( n558 )  ;
assign LB2D_proc_7_addr0 = n561 ? (LB2D_proc_x) : (0);
assign LB2D_proc_7_data0 = n561 ? (n217) : (LB2D_proc_7[0]);
function [7:0] gb_fun ;
input [647:0] arg0;
    begin
//TODO: Add the specific function HERE.    end
endfunction

always @(posedge clk) begin
   if(rst) begin
       LB1D_buff <= LB1D_buff;
       LB1D_p_cnt <= LB1D_p_cnt;
       LB2D_proc_w <= LB2D_proc_w;
       LB2D_proc_x <= LB2D_proc_x;
       LB2D_proc_y <= LB2D_proc_y;
       LB2D_shift_0 <= LB2D_shift_0;
       LB2D_shift_1 <= LB2D_shift_1;
       LB2D_shift_2 <= LB2D_shift_2;
       LB2D_shift_3 <= LB2D_shift_3;
       LB2D_shift_4 <= LB2D_shift_4;
       LB2D_shift_5 <= LB2D_shift_5;
       LB2D_shift_6 <= LB2D_shift_6;
       LB2D_shift_7 <= LB2D_shift_7;
       LB2D_shift_x <= LB2D_shift_x;
       LB2D_shift_y <= LB2D_shift_y;
       arg_0_TDATA <= arg_0_TDATA;
       arg_0_TVALID <= arg_0_TVALID;
       arg_1_TREADY <= arg_1_TREADY;
       gb_exit_it_1 <= gb_exit_it_1;
       gb_exit_it_2 <= gb_exit_it_2;
       gb_exit_it_3 <= gb_exit_it_3;
       gb_exit_it_4 <= gb_exit_it_4;
       gb_exit_it_5 <= gb_exit_it_5;
       gb_exit_it_6 <= gb_exit_it_6;
       gb_exit_it_7 <= gb_exit_it_7;
       gb_exit_it_8 <= gb_exit_it_8;
       gb_p_cnt <= gb_p_cnt;
       gb_pp_it_1 <= gb_pp_it_1;
       gb_pp_it_2 <= gb_pp_it_2;
       gb_pp_it_3 <= gb_pp_it_3;
       gb_pp_it_4 <= gb_pp_it_4;
       gb_pp_it_5 <= gb_pp_it_5;
       gb_pp_it_6 <= gb_pp_it_6;
       gb_pp_it_7 <= gb_pp_it_7;
       gb_pp_it_8 <= gb_pp_it_8;
       gb_pp_it_9 <= gb_pp_it_9;
       in_stream_buff_0 <= in_stream_buff_0;
       in_stream_buff_1 <= in_stream_buff_1;
       in_stream_empty <= in_stream_empty;
       in_stream_full <= in_stream_full;
       slice_stream_buff_0 <= slice_stream_buff_0;
       slice_stream_buff_1 <= slice_stream_buff_1;
       slice_stream_empty <= slice_stream_empty;
       slice_stream_full <= slice_stream_full;
       stencil_stream_buff_0 <= stencil_stream_buff_0;
       stencil_stream_buff_1 <= stencil_stream_buff_1;
       stencil_stream_empty <= stencil_stream_empty;
       stencil_stream_full <= stencil_stream_full;
   end
   else if(step) begin
       LB1D_buff <= n39;
       LB1D_p_cnt <= n41;
       LB2D_proc_w <= n52;
       LB2D_proc_x <= n60;
       LB2D_proc_y <= n70;
       LB2D_shift_0 <= n78;
       LB2D_shift_1 <= n84;
       LB2D_shift_2 <= n90;
       LB2D_shift_3 <= n96;
       LB2D_shift_4 <= n102;
       LB2D_shift_5 <= n108;
       LB2D_shift_6 <= n114;
       LB2D_shift_7 <= n120;
       LB2D_shift_x <= n129;
       LB2D_shift_y <= n139;
       arg_0_TDATA <= n148;
       arg_0_TVALID <= n156;
       arg_1_TREADY <= n165;
       gb_exit_it_1 <= n169;
       gb_exit_it_2 <= n170;
       gb_exit_it_3 <= n171;
       gb_exit_it_4 <= n172;
       gb_exit_it_5 <= n173;
       gb_exit_it_6 <= n174;
       gb_exit_it_7 <= n175;
       gb_exit_it_8 <= n176;
       gb_p_cnt <= n179;
       gb_pp_it_1 <= n180;
       gb_pp_it_2 <= n181;
       gb_pp_it_3 <= n182;
       gb_pp_it_4 <= n183;
       gb_pp_it_5 <= n184;
       gb_pp_it_6 <= n185;
       gb_pp_it_7 <= n186;
       gb_pp_it_8 <= n187;
       gb_pp_it_9 <= n188;
       in_stream_buff_0 <= n194;
       in_stream_buff_1 <= n200;
       in_stream_empty <= n208;
       in_stream_full <= n216;
       slice_stream_buff_0 <= n303;
       slice_stream_buff_1 <= n310;
       slice_stream_empty <= n318;
       slice_stream_full <= n327;
       stencil_stream_buff_0 <= n496;
       stencil_stream_buff_1 <= n502;
       stencil_stream_empty <= n510;
       stencil_stream_full <= n520;
       LB2D_proc_0 [ LB2D_proc_0_addr0 ] <= LB2D_proc_0_data0;
       LB2D_proc_1 [ LB2D_proc_1_addr0 ] <= LB2D_proc_1_data0;
       LB2D_proc_2 [ LB2D_proc_2_addr0 ] <= LB2D_proc_2_data0;
       LB2D_proc_3 [ LB2D_proc_3_addr0 ] <= LB2D_proc_3_data0;
       LB2D_proc_4 [ LB2D_proc_4_addr0 ] <= LB2D_proc_4_data0;
       LB2D_proc_5 [ LB2D_proc_5_addr0 ] <= LB2D_proc_5_data0;
       LB2D_proc_6 [ LB2D_proc_6_addr0 ] <= LB2D_proc_6_data0;
       LB2D_proc_7 [ LB2D_proc_7_addr0 ] <= LB2D_proc_7_data0;
   end
end
endmodule
