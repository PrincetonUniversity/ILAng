module alu(
pc,
r0,
r1,
r2,
r3,
clk,rst,
step
);
input clk;
input rst;
input step;
output      [7:0] pc;
output      [7:0] r0;
output      [7:0] r1;
output      [7:0] r2;
output      [7:0] r3;
reg      [7:0] pc;
reg      [7:0] r0;
reg      [7:0] r1;
reg      [7:0] r2;
reg      [7:0] r3;
wire      [7:0] n0;
wire      [5:0] n1;
wire            n2;
wire            n3;
wire            n4;
wire            n5;
wire            n6;
wire            n7;
wire            n8;
wire            n9;
wire            n10;
wire            n11;
wire            n12;
wire            n13;
wire            n14;
wire            n15;
wire            n16;
wire            n17;
wire            n18;
wire            n19;
wire            n20;
wire            n21;
wire            n22;
wire            n23;
wire            n24;
wire            n25;
wire            n26;
wire            n27;
wire            n28;
wire            n29;
wire            n30;
wire            n31;
wire            n32;
wire            n33;
wire            n34;
wire            n35;
wire            n36;
wire            n37;
wire            n38;
wire            n39;
wire            n40;
wire            n41;
wire            n42;
wire            n43;
wire            n44;
wire            n45;
wire            n46;
wire            n47;
wire            n48;
wire            n49;
wire            n50;
wire            n51;
wire            n52;
wire            n53;
wire            n54;
wire            n55;
wire            n56;
wire            n57;
wire            n58;
wire            n59;
wire            n60;
wire            n61;
wire            n62;
wire            n63;
wire            n64;
wire            n65;
wire            n66;
wire            n67;
wire            n68;
wire            n69;
wire            n70;
wire            n71;
wire            n72;
wire            n73;
wire            n74;
wire            n75;
wire            n76;
wire            n77;
wire            n78;
wire            n79;
wire            n80;
wire            n81;
wire            n82;
wire            n83;
wire            n84;
wire            n85;
wire            n86;
wire            n87;
wire            n88;
wire            n89;
wire            n90;
wire            n91;
wire            n92;
wire            n93;
wire            n94;
wire            n95;
wire            n96;
wire            n97;
wire            n98;
wire            n99;
wire            n100;
wire            n101;
wire            n102;
wire            n103;
wire            n104;
wire            n105;
wire            n106;
wire            n107;
wire            n108;
wire            n109;
wire            n110;
wire            n111;
wire            n112;
wire            n113;
wire            n114;
wire            n115;
wire            n116;
wire            n117;
wire            n118;
wire            n119;
wire            n120;
wire            n121;
wire            n122;
wire            n123;
wire            n124;
wire            n125;
wire            n126;
wire            n127;
wire            n128;
wire      [1:0] n129;
wire            n130;
wire            n131;
wire            n132;
wire      [7:0] n133;
wire      [7:0] n134;
wire      [7:0] n135;
wire      [7:0] n136;
wire            n137;
wire            n138;
wire            n139;
wire      [7:0] n140;
wire      [7:0] n141;
wire            n142;
wire            n143;
wire            n144;
wire      [7:0] n145;
wire      [7:0] n146;
wire      [7:0] n147;
wire      [7:0] n148;
wire      [7:0] n149;
wire      [7:0] n150;
wire      [7:0] n151;
wire      [7:0] n152;
wire      [7:0] n153;
wire      [7:0] n154;
wire      [7:0] n155;
wire      [7:0] n156;
wire      [7:0] n157;
wire      [7:0] n158;
wire      [7:0] n159;
wire      [7:0] n160;
wire      [7:0] n161;
wire      [7:0] n162;
wire      [7:0] n163;
wire            n164;
wire            n165;
wire            n166;
wire      [7:0] n167;
wire            n168;
wire            n169;
wire            n170;
wire      [7:0] n171;
wire      [7:0] n172;
wire      [7:0] n173;
wire      [7:0] n174;
wire      [7:0] n175;
wire      [7:0] n176;
wire      [7:0] n177;
wire      [7:0] n178;
wire      [7:0] n179;
wire      [7:0] n180;
wire      [7:0] n181;
wire      [7:0] n182;
wire      [7:0] n183;
wire      [7:0] n184;
wire      [7:0] n185;
wire      [7:0] n186;
wire      [7:0] n187;
wire      [7:0] n188;
wire            n189;
wire            n190;
wire            n191;
wire      [7:0] n192;
wire            n193;
wire            n194;
wire            n195;
wire      [7:0] n196;
wire      [7:0] n197;
wire      [7:0] n198;
wire      [7:0] n199;
wire      [7:0] n200;
wire      [7:0] n201;
wire      [7:0] n202;
wire      [7:0] n203;
wire      [7:0] n204;
wire      [7:0] n205;
wire      [7:0] n206;
wire      [7:0] n207;
wire      [7:0] n208;
wire      [7:0] n209;
wire      [7:0] n210;
wire      [7:0] n211;
wire            n212;
wire            n213;
wire            n214;
wire      [7:0] n215;
wire            n216;
wire            n217;
wire            n218;
wire      [7:0] n219;
wire      [7:0] n220;
wire      [7:0] n221;
wire      [7:0] n222;
wire      [7:0] n223;
wire      [7:0] n224;
wire      [7:0] n225;
wire      [7:0] n226;
wire      [7:0] n227;
wire      [7:0] n228;
wire      [7:0] n229;
wire      [7:0] n230;
wire      [7:0] n231;
wire      [7:0] n232;
wire      [7:0] n233;
wire      [7:0] n234;
wire      [7:0] n235;
reg      [7:0] rom[255:0];
wire clk;
wire rst;
wire step;
assign n0 =  (  rom [ pc ] )  ;
assign n1 = n0[5:0] ;
assign n2 =  ( n1 ) == ( 6'd63 )  ;
assign n3 =  ( n1 ) == ( 6'd62 )  ;
assign n4 =  ( n1 ) == ( 6'd61 )  ;
assign n5 =  ( n1 ) == ( 6'd60 )  ;
assign n6 =  ( n1 ) == ( 6'd59 )  ;
assign n7 =  ( n1 ) == ( 6'd58 )  ;
assign n8 =  ( n1 ) == ( 6'd57 )  ;
assign n9 =  ( n1 ) == ( 6'd56 )  ;
assign n10 =  ( n1 ) == ( 6'd55 )  ;
assign n11 =  ( n1 ) == ( 6'd54 )  ;
assign n12 =  ( n1 ) == ( 6'd53 )  ;
assign n13 =  ( n1 ) == ( 6'd52 )  ;
assign n14 =  ( n1 ) == ( 6'd51 )  ;
assign n15 =  ( n1 ) == ( 6'd50 )  ;
assign n16 =  ( n1 ) == ( 6'd49 )  ;
assign n17 =  ( n1 ) == ( 6'd48 )  ;
assign n18 =  ( n1 ) == ( 6'd47 )  ;
assign n19 =  ( n1 ) == ( 6'd46 )  ;
assign n20 =  ( n1 ) == ( 6'd45 )  ;
assign n21 =  ( n1 ) == ( 6'd44 )  ;
assign n22 =  ( n1 ) == ( 6'd43 )  ;
assign n23 =  ( n1 ) == ( 6'd42 )  ;
assign n24 =  ( n1 ) == ( 6'd41 )  ;
assign n25 =  ( n1 ) == ( 6'd40 )  ;
assign n26 =  ( n1 ) == ( 6'd39 )  ;
assign n27 =  ( n1 ) == ( 6'd38 )  ;
assign n28 =  ( n1 ) == ( 6'd37 )  ;
assign n29 =  ( n1 ) == ( 6'd36 )  ;
assign n30 =  ( n1 ) == ( 6'd35 )  ;
assign n31 =  ( n1 ) == ( 6'd34 )  ;
assign n32 =  ( n1 ) == ( 6'd33 )  ;
assign n33 =  ( n1 ) == ( 6'd32 )  ;
assign n34 =  ( n1 ) == ( 6'd31 )  ;
assign n35 =  ( n1 ) == ( 6'd30 )  ;
assign n36 =  ( n1 ) == ( 6'd29 )  ;
assign n37 =  ( n1 ) == ( 6'd28 )  ;
assign n38 =  ( n1 ) == ( 6'd27 )  ;
assign n39 =  ( n1 ) == ( 6'd26 )  ;
assign n40 =  ( n1 ) == ( 6'd25 )  ;
assign n41 =  ( n1 ) == ( 6'd24 )  ;
assign n42 =  ( n1 ) == ( 6'd23 )  ;
assign n43 =  ( n1 ) == ( 6'd22 )  ;
assign n44 =  ( n1 ) == ( 6'd21 )  ;
assign n45 =  ( n1 ) == ( 6'd20 )  ;
assign n46 =  ( n1 ) == ( 6'd19 )  ;
assign n47 =  ( n1 ) == ( 6'd18 )  ;
assign n48 =  ( n1 ) == ( 6'd17 )  ;
assign n49 =  ( n1 ) == ( 6'd16 )  ;
assign n50 =  ( n1 ) == ( 6'd15 )  ;
assign n51 =  ( n1 ) == ( 6'd14 )  ;
assign n52 =  ( n1 ) == ( 6'd13 )  ;
assign n53 =  ( n1 ) == ( 6'd12 )  ;
assign n54 =  ( n1 ) == ( 6'd11 )  ;
assign n55 =  ( n1 ) == ( 6'd10 )  ;
assign n56 =  ( n1 ) == ( 6'd9 )  ;
assign n57 =  ( n1 ) == ( 6'd8 )  ;
assign n58 =  ( n1 ) == ( 6'd7 )  ;
assign n59 =  ( n1 ) == ( 6'd6 )  ;
assign n60 =  ( n1 ) == ( 6'd5 )  ;
assign n61 =  ( n1 ) == ( 6'd4 )  ;
assign n62 =  ( n1 ) == ( 6'd3 )  ;
assign n63 =  ( n1 ) == ( 6'd2 )  ;
assign n64 =  ( n1 ) == ( 6'd1 )  ;
assign n65 =  ( n1 ) == ( 6'd0 )  ;
assign n66 =  ( n64 ) | ( n65 )  ;
assign n67 =  ( n63 ) | ( n66 )  ;
assign n68 =  ( n62 ) | ( n67 )  ;
assign n69 =  ( n61 ) | ( n68 )  ;
assign n70 =  ( n60 ) | ( n69 )  ;
assign n71 =  ( n59 ) | ( n70 )  ;
assign n72 =  ( n58 ) | ( n71 )  ;
assign n73 =  ( n57 ) | ( n72 )  ;
assign n74 =  ( n56 ) | ( n73 )  ;
assign n75 =  ( n55 ) | ( n74 )  ;
assign n76 =  ( n54 ) | ( n75 )  ;
assign n77 =  ( n53 ) | ( n76 )  ;
assign n78 =  ( n52 ) | ( n77 )  ;
assign n79 =  ( n51 ) | ( n78 )  ;
assign n80 =  ( n50 ) | ( n79 )  ;
assign n81 =  ( n49 ) | ( n80 )  ;
assign n82 =  ( n48 ) | ( n81 )  ;
assign n83 =  ( n47 ) | ( n82 )  ;
assign n84 =  ( n46 ) | ( n83 )  ;
assign n85 =  ( n45 ) | ( n84 )  ;
assign n86 =  ( n44 ) | ( n85 )  ;
assign n87 =  ( n43 ) | ( n86 )  ;
assign n88 =  ( n42 ) | ( n87 )  ;
assign n89 =  ( n41 ) | ( n88 )  ;
assign n90 =  ( n40 ) | ( n89 )  ;
assign n91 =  ( n39 ) | ( n90 )  ;
assign n92 =  ( n38 ) | ( n91 )  ;
assign n93 =  ( n37 ) | ( n92 )  ;
assign n94 =  ( n36 ) | ( n93 )  ;
assign n95 =  ( n35 ) | ( n94 )  ;
assign n96 =  ( n34 ) | ( n95 )  ;
assign n97 =  ( n33 ) | ( n96 )  ;
assign n98 =  ( n32 ) | ( n97 )  ;
assign n99 =  ( n31 ) | ( n98 )  ;
assign n100 =  ( n30 ) | ( n99 )  ;
assign n101 =  ( n29 ) | ( n100 )  ;
assign n102 =  ( n28 ) | ( n101 )  ;
assign n103 =  ( n27 ) | ( n102 )  ;
assign n104 =  ( n26 ) | ( n103 )  ;
assign n105 =  ( n25 ) | ( n104 )  ;
assign n106 =  ( n24 ) | ( n105 )  ;
assign n107 =  ( n23 ) | ( n106 )  ;
assign n108 =  ( n22 ) | ( n107 )  ;
assign n109 =  ( n21 ) | ( n108 )  ;
assign n110 =  ( n20 ) | ( n109 )  ;
assign n111 =  ( n19 ) | ( n110 )  ;
assign n112 =  ( n18 ) | ( n111 )  ;
assign n113 =  ( n17 ) | ( n112 )  ;
assign n114 =  ( n16 ) | ( n113 )  ;
assign n115 =  ( n15 ) | ( n114 )  ;
assign n116 =  ( n14 ) | ( n115 )  ;
assign n117 =  ( n13 ) | ( n116 )  ;
assign n118 =  ( n12 ) | ( n117 )  ;
assign n119 =  ( n11 ) | ( n118 )  ;
assign n120 =  ( n10 ) | ( n119 )  ;
assign n121 =  ( n9 ) | ( n120 )  ;
assign n122 =  ( n8 ) | ( n121 )  ;
assign n123 =  ( n7 ) | ( n122 )  ;
assign n124 =  ( n6 ) | ( n123 )  ;
assign n125 =  ( n5 ) | ( n124 )  ;
assign n126 =  ( n4 ) | ( n125 )  ;
assign n127 =  ( n3 ) | ( n126 )  ;
assign n128 =  ( n2 ) | ( n127 )  ;
assign n129 = n0[5:4] ;
assign n130 =  ( n129 ) == ( 2'd0 )  ;
assign n131 =  ( n129 ) == ( 2'd1 )  ;
assign n132 =  ( n130 ) | ( n131 )  ;
assign n133 =  ( pc ) + ( 8'd1 )  ;
assign n134 =  ( pc ) + ( 8'd2 )  ;
assign n135 =  ( n132 ) ? ( n133 ) : ( n134 ) ;
assign n136 =  ( n128 ) ? ( n135 ) : ( pc ) ;
assign n137 =  ( n13 ) | ( n17 )  ;
assign n138 =  ( n9 ) | ( n137 )  ;
assign n139 =  ( n5 ) | ( n138 )  ;
assign n140 =  (  rom [ n133 ] )  ;
assign n141 =  ( r0 ) - ( n140 )  ;
assign n142 =  ( n29 ) | ( n33 )  ;
assign n143 =  ( n25 ) | ( n142 )  ;
assign n144 =  ( n21 ) | ( n143 )  ;
assign n145 =  ( r0 ) + ( n140 )  ;
assign n146 =  ( r0 ) - ( r3 )  ;
assign n147 =  ( r0 ) - ( r2 )  ;
assign n148 =  ( r0 ) - ( r1 )  ;
assign n149 =  ( r3 ) - ( r3 )  ;
assign n150 =  ( r3 ) + ( r0 )  ;
assign n151 =  ( r0 ) + ( r2 )  ;
assign n152 =  ( r0 ) + ( r1 )  ;
assign n153 =  ( r0 ) + ( r0 )  ;
assign n154 =  ( n65 ) ? ( n153 ) : ( r0 ) ;
assign n155 =  ( n61 ) ? ( n152 ) : ( n154 ) ;
assign n156 =  ( n57 ) ? ( n151 ) : ( n155 ) ;
assign n157 =  ( n53 ) ? ( n150 ) : ( n156 ) ;
assign n158 =  ( n49 ) ? ( n149 ) : ( n157 ) ;
assign n159 =  ( n45 ) ? ( n148 ) : ( n158 ) ;
assign n160 =  ( n41 ) ? ( n147 ) : ( n159 ) ;
assign n161 =  ( n37 ) ? ( n146 ) : ( n160 ) ;
assign n162 =  ( n144 ) ? ( n145 ) : ( n161 ) ;
assign n163 =  ( n139 ) ? ( n141 ) : ( n162 ) ;
assign n164 =  ( n12 ) | ( n16 )  ;
assign n165 =  ( n8 ) | ( n164 )  ;
assign n166 =  ( n4 ) | ( n165 )  ;
assign n167 =  ( r1 ) - ( n140 )  ;
assign n168 =  ( n28 ) | ( n32 )  ;
assign n169 =  ( n24 ) | ( n168 )  ;
assign n170 =  ( n20 ) | ( n169 )  ;
assign n171 =  ( r1 ) + ( n140 )  ;
assign n172 =  ( r1 ) - ( r3 )  ;
assign n173 =  ( r1 ) - ( r2 )  ;
assign n174 =  ( r1 ) - ( r0 )  ;
assign n175 =  ( r3 ) + ( r1 )  ;
assign n176 =  ( r2 ) + ( r1 )  ;
assign n177 =  ( r1 ) + ( r1 )  ;
assign n178 =  ( r1 ) + ( r0 )  ;
assign n179 =  ( n64 ) ? ( n178 ) : ( r1 ) ;
assign n180 =  ( n60 ) ? ( n177 ) : ( n179 ) ;
assign n181 =  ( n56 ) ? ( n176 ) : ( n180 ) ;
assign n182 =  ( n52 ) ? ( n175 ) : ( n181 ) ;
assign n183 =  ( n48 ) ? ( n174 ) : ( n182 ) ;
assign n184 =  ( n44 ) ? ( n149 ) : ( n183 ) ;
assign n185 =  ( n40 ) ? ( n173 ) : ( n184 ) ;
assign n186 =  ( n36 ) ? ( n172 ) : ( n185 ) ;
assign n187 =  ( n170 ) ? ( n171 ) : ( n186 ) ;
assign n188 =  ( n166 ) ? ( n167 ) : ( n187 ) ;
assign n189 =  ( n11 ) | ( n15 )  ;
assign n190 =  ( n7 ) | ( n189 )  ;
assign n191 =  ( n3 ) | ( n190 )  ;
assign n192 =  ( r2 ) - ( n140 )  ;
assign n193 =  ( n27 ) | ( n31 )  ;
assign n194 =  ( n23 ) | ( n193 )  ;
assign n195 =  ( n19 ) | ( n194 )  ;
assign n196 =  ( r2 ) + ( n140 )  ;
assign n197 =  ( r2 ) - ( r3 )  ;
assign n198 =  ( r2 ) - ( r1 )  ;
assign n199 =  ( r2 ) - ( r0 )  ;
assign n200 =  ( r3 ) + ( r2 )  ;
assign n201 =  ( r2 ) + ( r2 )  ;
assign n202 =  ( n63 ) ? ( n151 ) : ( r2 ) ;
assign n203 =  ( n59 ) ? ( n176 ) : ( n202 ) ;
assign n204 =  ( n55 ) ? ( n201 ) : ( n203 ) ;
assign n205 =  ( n51 ) ? ( n200 ) : ( n204 ) ;
assign n206 =  ( n47 ) ? ( n199 ) : ( n205 ) ;
assign n207 =  ( n43 ) ? ( n198 ) : ( n206 ) ;
assign n208 =  ( n39 ) ? ( n149 ) : ( n207 ) ;
assign n209 =  ( n35 ) ? ( n197 ) : ( n208 ) ;
assign n210 =  ( n195 ) ? ( n196 ) : ( n209 ) ;
assign n211 =  ( n191 ) ? ( n192 ) : ( n210 ) ;
assign n212 =  ( n10 ) | ( n14 )  ;
assign n213 =  ( n6 ) | ( n212 )  ;
assign n214 =  ( n2 ) | ( n213 )  ;
assign n215 =  ( r3 ) - ( n140 )  ;
assign n216 =  ( n26 ) | ( n30 )  ;
assign n217 =  ( n22 ) | ( n216 )  ;
assign n218 =  ( n18 ) | ( n217 )  ;
assign n219 =  ( r3 ) + ( n140 )  ;
assign n220 =  ( r3 ) - ( r2 )  ;
assign n221 =  ( r3 ) - ( r1 )  ;
assign n222 =  ( r3 ) - ( r0 )  ;
assign n223 =  ( r3 ) + ( r3 )  ;
assign n224 =  ( r1 ) + ( r3 )  ;
assign n225 =  ( r0 ) + ( r3 )  ;
assign n226 =  ( n62 ) ? ( n225 ) : ( r3 ) ;
assign n227 =  ( n58 ) ? ( n224 ) : ( n226 ) ;
assign n228 =  ( n54 ) ? ( n200 ) : ( n227 ) ;
assign n229 =  ( n50 ) ? ( n223 ) : ( n228 ) ;
assign n230 =  ( n46 ) ? ( n222 ) : ( n229 ) ;
assign n231 =  ( n42 ) ? ( n221 ) : ( n230 ) ;
assign n232 =  ( n38 ) ? ( n220 ) : ( n231 ) ;
assign n233 =  ( n34 ) ? ( n149 ) : ( n232 ) ;
assign n234 =  ( n218 ) ? ( n219 ) : ( n233 ) ;
assign n235 =  ( n214 ) ? ( n215 ) : ( n234 ) ;
always @(posedge clk) begin
   if(rst) begin
       pc <= pc;
       r0 <= r0;
       r1 <= r1;
       r2 <= r2;
       r3 <= r3;
   end
   else if(step) begin
       pc <= n136;
       r0 <= n163;
       r1 <= n188;
       r2 <= n211;
       r3 <= n235;
   end
end
endmodule
