module GB(
arg_0_TREADY,
arg_1_TDATA,
arg_1_TVALID,
LB1D_buff,
LB1D_in,
LB1D_it_1,
LB1D_p_cnt,
LB2D_proc_w,
LB2D_proc_x,
LB2D_proc_y,
LB2D_shift_0,
LB2D_shift_1,
LB2D_shift_2,
LB2D_shift_3,
LB2D_shift_4,
LB2D_shift_5,
LB2D_shift_6,
LB2D_shift_7,
LB2D_shift_x,
LB2D_shift_y,
arg_0_TDATA,
arg_0_TVALID,
arg_1_TREADY,
gb_exit_it_1,
gb_exit_it_2,
gb_exit_it_3,
gb_exit_it_4,
gb_exit_it_5,
gb_exit_it_6,
gb_exit_it_7,
gb_exit_it_8,
gb_p_cnt,
gb_pp_it_1,
gb_pp_it_2,
gb_pp_it_3,
gb_pp_it_4,
gb_pp_it_5,
gb_pp_it_6,
gb_pp_it_7,
gb_pp_it_8,
gb_pp_it_9,
in_stream_buff_0,
in_stream_buff_1,
in_stream_empty,
in_stream_full,
slice_stream_buff_0,
slice_stream_buff_1,
slice_stream_empty,
slice_stream_full,
stencil_stream_buff_0,
stencil_stream_buff_1,
stencil_stream_empty,
stencil_stream_full,
clk,rst,
step
);
input            arg_0_TREADY;
input      [7:0] arg_1_TDATA;
input            arg_1_TVALID;
input clk;
input rst;
input step;
output      [7:0] LB1D_buff;
output      [7:0] LB1D_in;
output            LB1D_it_1;
output     [18:0] LB1D_p_cnt;
output     [63:0] LB2D_proc_w;
output      [8:0] LB2D_proc_x;
output      [9:0] LB2D_proc_y;
output     [71:0] LB2D_shift_0;
output     [71:0] LB2D_shift_1;
output     [71:0] LB2D_shift_2;
output     [71:0] LB2D_shift_3;
output     [71:0] LB2D_shift_4;
output     [71:0] LB2D_shift_5;
output     [71:0] LB2D_shift_6;
output     [71:0] LB2D_shift_7;
output      [8:0] LB2D_shift_x;
output      [9:0] LB2D_shift_y;
output      [7:0] arg_0_TDATA;
output            arg_0_TVALID;
output            arg_1_TREADY;
output            gb_exit_it_1;
output            gb_exit_it_2;
output            gb_exit_it_3;
output            gb_exit_it_4;
output            gb_exit_it_5;
output            gb_exit_it_6;
output            gb_exit_it_7;
output            gb_exit_it_8;
output     [18:0] gb_p_cnt;
output            gb_pp_it_1;
output            gb_pp_it_2;
output            gb_pp_it_3;
output            gb_pp_it_4;
output            gb_pp_it_5;
output            gb_pp_it_6;
output            gb_pp_it_7;
output            gb_pp_it_8;
output            gb_pp_it_9;
output      [7:0] in_stream_buff_0;
output      [7:0] in_stream_buff_1;
output            in_stream_empty;
output            in_stream_full;
output     [71:0] slice_stream_buff_0;
output     [71:0] slice_stream_buff_1;
output            slice_stream_empty;
output            slice_stream_full;
output    [647:0] stencil_stream_buff_0;
output    [647:0] stencil_stream_buff_1;
output            stencil_stream_empty;
output            stencil_stream_full;
reg      [7:0] LB1D_buff;
reg      [7:0] LB1D_in;
reg            LB1D_it_1;
reg     [18:0] LB1D_p_cnt;
reg     [63:0] LB2D_proc_w;
reg      [8:0] LB2D_proc_x;
reg      [9:0] LB2D_proc_y;
reg     [71:0] LB2D_shift_0;
reg     [71:0] LB2D_shift_1;
reg     [71:0] LB2D_shift_2;
reg     [71:0] LB2D_shift_3;
reg     [71:0] LB2D_shift_4;
reg     [71:0] LB2D_shift_5;
reg     [71:0] LB2D_shift_6;
reg     [71:0] LB2D_shift_7;
reg      [8:0] LB2D_shift_x;
reg      [9:0] LB2D_shift_y;
reg      [7:0] arg_0_TDATA;
reg            arg_0_TVALID;
reg            arg_1_TREADY;
reg            gb_exit_it_1;
reg            gb_exit_it_2;
reg            gb_exit_it_3;
reg            gb_exit_it_4;
reg            gb_exit_it_5;
reg            gb_exit_it_6;
reg            gb_exit_it_7;
reg            gb_exit_it_8;
reg     [18:0] gb_p_cnt;
reg            gb_pp_it_1;
reg            gb_pp_it_2;
reg            gb_pp_it_3;
reg            gb_pp_it_4;
reg            gb_pp_it_5;
reg            gb_pp_it_6;
reg            gb_pp_it_7;
reg            gb_pp_it_8;
reg            gb_pp_it_9;
reg      [7:0] in_stream_buff_0;
reg      [7:0] in_stream_buff_1;
reg            in_stream_empty;
reg            in_stream_full;
reg     [71:0] slice_stream_buff_0;
reg     [71:0] slice_stream_buff_1;
reg            slice_stream_empty;
reg            slice_stream_full;
reg    [647:0] stencil_stream_buff_0;
reg    [647:0] stencil_stream_buff_1;
reg            stencil_stream_empty;
reg            stencil_stream_full;
wire            arg_0_TREADY;
wire      [7:0] arg_1_TDATA;
wire            arg_1_TVALID;
wire            n0;
wire            n1;
wire            n2;
wire            n3;
wire            n4;
wire            n5;
wire            n6;
wire            n7;
wire            n8;
wire            n9;
wire            n10;
wire            n11;
wire            n12;
wire            n13;
wire            n14;
wire            n15;
wire            n16;
wire            n17;
wire            n18;
wire            n19;
wire            n20;
wire            n21;
wire            n22;
wire            n23;
wire            n24;
wire            n25;
wire            n26;
wire            n27;
wire            n28;
wire            n29;
wire            n30;
wire            n31;
wire            n32;
wire            n33;
wire            n34;
wire            n35;
wire            n36;
wire            n37;
wire      [7:0] n38;
wire      [7:0] n39;
wire      [7:0] n40;
wire      [7:0] n41;
wire      [7:0] n42;
wire      [7:0] n43;
wire      [7:0] n44;
wire      [7:0] n45;
wire      [7:0] n46;
wire      [7:0] n47;
wire      [7:0] n48;
wire      [7:0] n49;
wire            n50;
wire            n51;
wire            n52;
wire     [18:0] n53;
wire     [18:0] n54;
wire            n55;
wire     [18:0] n56;
wire     [18:0] n57;
wire     [18:0] n58;
wire     [18:0] n59;
wire     [18:0] n60;
wire     [18:0] n61;
wire     [18:0] n62;
wire     [18:0] n63;
wire            n64;
wire            n65;
wire     [63:0] n66;
wire     [63:0] n67;
wire     [63:0] n68;
wire     [63:0] n69;
wire     [63:0] n70;
wire     [63:0] n71;
wire     [63:0] n72;
wire     [63:0] n73;
wire     [63:0] n74;
wire            n75;
wire            n76;
wire            n77;
wire      [8:0] n78;
wire      [8:0] n79;
wire      [8:0] n80;
wire      [8:0] n81;
wire      [8:0] n82;
wire      [8:0] n83;
wire      [8:0] n84;
wire      [8:0] n85;
wire            n86;
wire      [9:0] n87;
wire      [9:0] n88;
wire      [9:0] n89;
wire      [9:0] n90;
wire      [9:0] n91;
wire      [9:0] n92;
wire      [9:0] n93;
wire            n94;
wire     [71:0] n95;
wire     [71:0] n96;
wire     [71:0] n97;
wire     [71:0] n98;
wire     [71:0] n99;
wire     [71:0] n100;
wire     [71:0] n101;
wire     [71:0] n102;
wire     [71:0] n103;
wire     [71:0] n104;
wire     [71:0] n105;
wire     [71:0] n106;
wire     [71:0] n107;
wire     [71:0] n108;
wire     [71:0] n109;
wire     [71:0] n110;
wire     [71:0] n111;
wire     [71:0] n112;
wire     [71:0] n113;
wire     [71:0] n114;
wire     [71:0] n115;
wire     [71:0] n116;
wire     [71:0] n117;
wire     [71:0] n118;
wire     [71:0] n119;
wire     [71:0] n120;
wire     [71:0] n121;
wire     [71:0] n122;
wire     [71:0] n123;
wire     [71:0] n124;
wire     [71:0] n125;
wire     [71:0] n126;
wire     [71:0] n127;
wire     [71:0] n128;
wire     [71:0] n129;
wire     [71:0] n130;
wire     [71:0] n131;
wire     [71:0] n132;
wire     [71:0] n133;
wire     [71:0] n134;
wire     [71:0] n135;
wire     [71:0] n136;
wire     [71:0] n137;
wire     [71:0] n138;
wire     [71:0] n139;
wire     [71:0] n140;
wire     [71:0] n141;
wire     [71:0] n142;
wire     [71:0] n143;
wire      [8:0] n144;
wire      [8:0] n145;
wire      [8:0] n146;
wire      [8:0] n147;
wire      [8:0] n148;
wire      [8:0] n149;
wire      [8:0] n150;
wire            n151;
wire            n152;
wire      [9:0] n153;
wire      [9:0] n154;
wire      [9:0] n155;
wire      [9:0] n156;
wire      [9:0] n157;
wire      [9:0] n158;
wire      [9:0] n159;
wire      [9:0] n160;
wire      [9:0] n161;
wire            n162;
wire    [647:0] n163;
wire      [7:0] n164;
wire      [7:0] n165;
wire      [7:0] n166;
wire      [7:0] n167;
wire      [7:0] n168;
wire      [7:0] n169;
wire      [7:0] n170;
wire            n171;
wire            n172;
wire            n173;
wire            n174;
wire            n175;
wire            n176;
wire            n177;
wire            n178;
wire            n179;
wire            n180;
wire            n181;
wire            n182;
wire            n183;
wire            n184;
wire            n185;
wire     [18:0] n186;
wire            n187;
wire            n188;
wire            n189;
wire            n190;
wire            n191;
wire            n192;
wire            n193;
wire            n194;
wire            n195;
wire            n196;
wire            n197;
wire            n198;
wire            n199;
wire            n200;
wire            n201;
wire            n202;
wire            n203;
wire            n204;
wire            n205;
wire            n206;
wire            n207;
wire            n208;
wire            n209;
wire            n210;
wire            n211;
wire            n212;
wire            n213;
wire            n214;
wire            n215;
wire            n216;
wire            n217;
wire            n218;
wire            n219;
wire            n220;
wire            n221;
wire            n222;
wire            n223;
wire            n224;
wire            n225;
wire            n226;
wire            n227;
wire            n228;
wire            n229;
wire            n230;
wire            n231;
wire            n232;
wire            n233;
wire            n234;
wire            n235;
wire            n236;
wire            n237;
wire     [18:0] n238;
wire     [18:0] n239;
wire     [18:0] n240;
wire     [18:0] n241;
wire     [18:0] n242;
wire     [18:0] n243;
wire     [18:0] n244;
wire            n245;
wire            n246;
wire            n247;
wire            n248;
wire            n249;
wire            n250;
wire            n251;
wire            n252;
wire            n253;
wire            n254;
wire            n255;
wire            n256;
wire            n257;
wire            n258;
wire            n259;
wire            n260;
wire            n261;
wire            n262;
wire            n263;
wire            n264;
wire            n265;
wire            n266;
wire            n267;
wire            n268;
wire            n269;
wire            n270;
wire            n271;
wire            n272;
wire            n273;
wire            n274;
wire            n275;
wire            n276;
wire            n277;
wire            n278;
wire            n279;
wire            n280;
wire            n281;
wire            n282;
wire            n283;
wire            n284;
wire            n285;
wire            n286;
wire            n287;
wire            n288;
wire            n289;
wire            n290;
wire            n291;
wire            n292;
wire            n293;
wire            n294;
wire            n295;
wire            n296;
wire            n297;
wire            n298;
wire      [7:0] n299;
wire      [7:0] n300;
wire      [7:0] n301;
wire      [7:0] n302;
wire      [7:0] n303;
wire      [7:0] n304;
wire      [7:0] n305;
wire      [7:0] n306;
wire      [7:0] n307;
wire      [7:0] n308;
wire      [7:0] n309;
wire      [7:0] n310;
wire            n311;
wire            n312;
wire            n313;
wire            n314;
wire            n315;
wire            n316;
wire            n317;
wire            n318;
wire            n319;
wire            n320;
wire            n321;
wire            n322;
wire            n323;
wire            n324;
wire            n325;
wire            n326;
wire      [7:0] n327;
wire            n328;
wire      [7:0] n329;
wire            n330;
wire      [7:0] n331;
wire            n332;
wire      [7:0] n333;
wire            n334;
wire      [7:0] n335;
wire            n336;
wire      [7:0] n337;
wire            n338;
wire      [7:0] n339;
wire            n340;
wire      [7:0] n341;
wire      [7:0] n342;
wire      [7:0] n343;
wire      [7:0] n344;
wire      [7:0] n345;
wire      [7:0] n346;
wire      [7:0] n347;
wire      [7:0] n348;
wire      [7:0] n349;
wire      [7:0] n350;
wire      [7:0] n351;
wire      [7:0] n352;
wire      [7:0] n353;
wire      [7:0] n354;
wire      [7:0] n355;
wire      [7:0] n356;
wire      [7:0] n357;
wire      [7:0] n358;
wire      [7:0] n359;
wire      [7:0] n360;
wire      [7:0] n361;
wire      [7:0] n362;
wire      [7:0] n363;
wire      [7:0] n364;
wire      [7:0] n365;
wire      [7:0] n366;
wire      [7:0] n367;
wire      [7:0] n368;
wire      [7:0] n369;
wire      [7:0] n370;
wire      [7:0] n371;
wire      [7:0] n372;
wire      [7:0] n373;
wire      [7:0] n374;
wire      [7:0] n375;
wire      [7:0] n376;
wire      [7:0] n377;
wire      [7:0] n378;
wire      [7:0] n379;
wire      [7:0] n380;
wire      [7:0] n381;
wire      [7:0] n382;
wire      [7:0] n383;
wire      [7:0] n384;
wire      [7:0] n385;
wire      [7:0] n386;
wire      [7:0] n387;
wire      [7:0] n388;
wire      [7:0] n389;
wire      [7:0] n390;
wire      [7:0] n391;
wire      [7:0] n392;
wire      [7:0] n393;
wire      [7:0] n394;
wire      [7:0] n395;
wire      [7:0] n396;
wire      [7:0] n397;
wire      [7:0] n398;
wire     [15:0] n399;
wire     [23:0] n400;
wire     [31:0] n401;
wire     [39:0] n402;
wire     [47:0] n403;
wire     [55:0] n404;
wire     [63:0] n405;
wire     [71:0] n406;
wire     [71:0] n407;
wire     [71:0] n408;
wire     [71:0] n409;
wire     [71:0] n410;
wire     [71:0] n411;
wire     [71:0] n412;
wire     [71:0] n413;
wire     [71:0] n414;
wire     [71:0] n415;
wire     [71:0] n416;
wire     [71:0] n417;
wire     [71:0] n418;
wire     [71:0] n419;
wire     [71:0] n420;
wire            n421;
wire            n422;
wire            n423;
wire            n424;
wire            n425;
wire            n426;
wire            n427;
wire            n428;
wire            n429;
wire            n430;
wire            n431;
wire            n432;
wire            n433;
wire            n434;
wire            n435;
wire            n436;
wire            n437;
wire            n438;
wire      [7:0] n439;
wire      [7:0] n440;
wire      [7:0] n441;
wire      [7:0] n442;
wire      [7:0] n443;
wire      [7:0] n444;
wire      [7:0] n445;
wire      [7:0] n446;
wire      [7:0] n447;
wire     [15:0] n448;
wire     [23:0] n449;
wire     [31:0] n450;
wire     [39:0] n451;
wire     [47:0] n452;
wire     [55:0] n453;
wire     [63:0] n454;
wire     [71:0] n455;
wire      [7:0] n456;
wire      [7:0] n457;
wire      [7:0] n458;
wire      [7:0] n459;
wire      [7:0] n460;
wire      [7:0] n461;
wire      [7:0] n462;
wire      [7:0] n463;
wire      [7:0] n464;
wire     [15:0] n465;
wire     [23:0] n466;
wire     [31:0] n467;
wire     [39:0] n468;
wire     [47:0] n469;
wire     [55:0] n470;
wire     [63:0] n471;
wire     [71:0] n472;
wire      [7:0] n473;
wire      [7:0] n474;
wire      [7:0] n475;
wire      [7:0] n476;
wire      [7:0] n477;
wire      [7:0] n478;
wire      [7:0] n479;
wire      [7:0] n480;
wire      [7:0] n481;
wire     [15:0] n482;
wire     [23:0] n483;
wire     [31:0] n484;
wire     [39:0] n485;
wire     [47:0] n486;
wire     [55:0] n487;
wire     [63:0] n488;
wire     [71:0] n489;
wire      [7:0] n490;
wire      [7:0] n491;
wire      [7:0] n492;
wire      [7:0] n493;
wire      [7:0] n494;
wire      [7:0] n495;
wire      [7:0] n496;
wire      [7:0] n497;
wire      [7:0] n498;
wire     [15:0] n499;
wire     [23:0] n500;
wire     [31:0] n501;
wire     [39:0] n502;
wire     [47:0] n503;
wire     [55:0] n504;
wire     [63:0] n505;
wire     [71:0] n506;
wire      [7:0] n507;
wire      [7:0] n508;
wire      [7:0] n509;
wire      [7:0] n510;
wire      [7:0] n511;
wire      [7:0] n512;
wire      [7:0] n513;
wire      [7:0] n514;
wire      [7:0] n515;
wire     [15:0] n516;
wire     [23:0] n517;
wire     [31:0] n518;
wire     [39:0] n519;
wire     [47:0] n520;
wire     [55:0] n521;
wire     [63:0] n522;
wire     [71:0] n523;
wire      [7:0] n524;
wire      [7:0] n525;
wire      [7:0] n526;
wire      [7:0] n527;
wire      [7:0] n528;
wire      [7:0] n529;
wire      [7:0] n530;
wire      [7:0] n531;
wire      [7:0] n532;
wire     [15:0] n533;
wire     [23:0] n534;
wire     [31:0] n535;
wire     [39:0] n536;
wire     [47:0] n537;
wire     [55:0] n538;
wire     [63:0] n539;
wire     [71:0] n540;
wire      [7:0] n541;
wire      [7:0] n542;
wire      [7:0] n543;
wire      [7:0] n544;
wire      [7:0] n545;
wire      [7:0] n546;
wire      [7:0] n547;
wire      [7:0] n548;
wire      [7:0] n549;
wire     [15:0] n550;
wire     [23:0] n551;
wire     [31:0] n552;
wire     [39:0] n553;
wire     [47:0] n554;
wire     [55:0] n555;
wire     [63:0] n556;
wire     [71:0] n557;
wire      [7:0] n558;
wire      [7:0] n559;
wire      [7:0] n560;
wire      [7:0] n561;
wire      [7:0] n562;
wire      [7:0] n563;
wire      [7:0] n564;
wire      [7:0] n565;
wire      [7:0] n566;
wire     [15:0] n567;
wire     [23:0] n568;
wire     [31:0] n569;
wire     [39:0] n570;
wire     [47:0] n571;
wire     [55:0] n572;
wire     [63:0] n573;
wire     [71:0] n574;
wire      [7:0] n575;
wire      [7:0] n576;
wire      [7:0] n577;
wire      [7:0] n578;
wire      [7:0] n579;
wire      [7:0] n580;
wire      [7:0] n581;
wire      [7:0] n582;
wire      [7:0] n583;
wire     [15:0] n584;
wire     [23:0] n585;
wire     [31:0] n586;
wire     [39:0] n587;
wire     [47:0] n588;
wire     [55:0] n589;
wire     [63:0] n590;
wire     [71:0] n591;
wire    [143:0] n592;
wire    [215:0] n593;
wire    [287:0] n594;
wire    [359:0] n595;
wire    [431:0] n596;
wire    [503:0] n597;
wire    [575:0] n598;
wire    [647:0] n599;
wire    [647:0] n600;
wire    [647:0] n601;
wire    [647:0] n602;
wire    [647:0] n603;
wire    [647:0] n604;
wire    [647:0] n605;
wire    [647:0] n606;
wire    [647:0] n607;
wire    [647:0] n608;
wire    [647:0] n609;
wire    [647:0] n610;
wire    [647:0] n611;
wire    [647:0] n612;
wire            n613;
wire            n614;
wire            n615;
wire            n616;
wire            n617;
wire            n618;
wire            n619;
wire            n620;
wire            n621;
wire            n622;
wire            n623;
wire            n624;
wire            n625;
wire            n626;
wire            n627;
wire            n628;
wire            n629;
wire            n630;
wire      [8:0] LB2D_proc_0_addr0;
wire      [7:0] LB2D_proc_0_data0;
wire            n631;
wire            n632;
wire            n633;
wire            n634;
wire            n635;
wire            n636;
wire            n637;
wire            n638;
wire            n639;
wire            n640;
wire            n641;
wire            n642;
wire            n643;
wire            n644;
wire            n645;
wire            n646;
wire            n647;
wire            n648;
wire            n649;
wire      [8:0] LB2D_proc_1_addr0;
wire      [7:0] LB2D_proc_1_data0;
wire            n650;
wire            n651;
wire            n652;
wire      [8:0] LB2D_proc_2_addr0;
wire      [7:0] LB2D_proc_2_data0;
wire            n653;
wire            n654;
wire            n655;
wire      [8:0] LB2D_proc_3_addr0;
wire      [7:0] LB2D_proc_3_data0;
wire            n656;
wire            n657;
wire            n658;
wire      [8:0] LB2D_proc_4_addr0;
wire      [7:0] LB2D_proc_4_data0;
wire            n659;
wire            n660;
wire            n661;
wire      [8:0] LB2D_proc_5_addr0;
wire      [7:0] LB2D_proc_5_data0;
wire            n662;
wire            n663;
wire            n664;
wire      [8:0] LB2D_proc_6_addr0;
wire      [7:0] LB2D_proc_6_data0;
wire            n665;
wire            n666;
wire            n667;
wire      [8:0] LB2D_proc_7_addr0;
wire      [7:0] LB2D_proc_7_data0;
wire            n668;
wire            n669;
wire            n670;
wire            n671;
reg      [7:0] LB2D_proc_0[511:0];
reg      [7:0] LB2D_proc_1[511:0];
reg      [7:0] LB2D_proc_2[511:0];
reg      [7:0] LB2D_proc_3[511:0];
reg      [7:0] LB2D_proc_4[511:0];
reg      [7:0] LB2D_proc_5[511:0];
reg      [7:0] LB2D_proc_6[511:0];
reg      [7:0] LB2D_proc_7[511:0];
wire clk;
wire rst;
wire step;
assign n0 =  ( arg_0_TREADY ) == ( 1'd1 )  ;
assign n1 =  ( arg_0_TVALID ) == ( 1'd1 )  ;
assign n2 =  ( n0 ) & ( n1 )  ;
assign n3 =  ( arg_1_TVALID ) == ( 1'd0 )  ;
assign n4 =  ( n2 ) & ( n3 )  ;
assign n5 =  ( arg_1_TREADY ) == ( 1'd1 )  ;
assign n6 =  ( arg_1_TVALID ) == ( 1'd1 )  ;
assign n7 =  ( n5 ) & ( n6 )  ;
assign n8 =  ( arg_0_TREADY ) == ( 1'd0 )  ;
assign n9 =  ( n7 ) & ( n8 )  ;
assign n10 =  ( arg_0_TVALID ) == ( 1'd0 )  ;
assign n11 =  ( gb_exit_it_1 ) == ( 1'd0 )  ;
assign n12 =  ( stencil_stream_empty ) == ( 1'd0 )  ;
assign n13 =  ( n11 ) & ( n12 )  ;
assign n14 =  ( gb_exit_it_1 ) == ( 1'd1 )  ;
assign n15 =  ( gb_exit_it_8 ) == ( 1'd0 )  ;
assign n16 =  ( n14 ) & ( n15 )  ;
assign n17 =  ( n13 ) | ( n16 )  ;
assign n18 =  ( n10 ) & ( n17 )  ;
assign n19 =  ( slice_stream_empty ) == ( 1'd0 )  ;
assign n20 =  ( LB2D_shift_x ) != ( 9'd488 )  ;
assign n21 =  ( n19 ) & ( n20 )  ;
assign n22 =  ( stencil_stream_full ) == ( 1'd0 )  ;
assign n23 =  ( LB2D_shift_x ) < ( 9'd8 )  ;
assign n24 =  ( n22 ) | ( n23 )  ;
assign n25 =  ( n21 ) & ( n24 )  ;
assign n26 =  ( in_stream_empty ) == ( 1'd0 )  ;
assign n27 =  ( LB2D_proc_x ) != ( 9'd488 )  ;
assign n28 =  ( n26 ) & ( n27 )  ;
assign n29 =  ( slice_stream_full ) == ( 1'd0 )  ;
assign n30 =  ( LB2D_proc_y ) < ( 10'd8 )  ;
assign n31 =  ( n29 ) | ( n30 )  ;
assign n32 =  ( n28 ) & ( n31 )  ;
assign n33 =  ( arg_1_TREADY ) == ( 1'd0 )  ;
assign n34 =  ( in_stream_full ) == ( 1'd0 )  ;
assign n35 =  ( n33 ) & ( n34 )  ;
assign n36 =  ( LB1D_it_1 ) == ( 1'd1 )  ;
assign n37 =  ( n35 ) & ( n36 )  ;
assign n38 =  ( n37 ) ? ( LB1D_in ) : ( LB1D_buff ) ;
assign n39 =  ( n32 ) ? ( LB1D_buff ) : ( n38 ) ;
assign n40 =  ( n25 ) ? ( LB1D_buff ) : ( n39 ) ;
assign n41 =  ( n18 ) ? ( LB1D_buff ) : ( n40 ) ;
assign n42 =  ( n9 ) ? ( LB1D_buff ) : ( n41 ) ;
assign n43 =  ( n4 ) ? ( LB1D_buff ) : ( n42 ) ;
assign n44 =  ( n37 ) ? ( arg_1_TDATA ) : ( LB1D_in ) ;
assign n45 =  ( n32 ) ? ( LB1D_in ) : ( n44 ) ;
assign n46 =  ( n25 ) ? ( LB1D_in ) : ( n45 ) ;
assign n47 =  ( n18 ) ? ( LB1D_in ) : ( n46 ) ;
assign n48 =  ( n9 ) ? ( LB1D_in ) : ( n47 ) ;
assign n49 =  ( n4 ) ? ( LB1D_in ) : ( n48 ) ;
assign n50 =  ( LB1D_it_1 ) == ( 1'd0 )  ;
assign n51 =  ( n35 ) & ( n50 )  ;
assign n52 =  ( n51 ) ? ( 1'd1 ) : ( LB1D_it_1 ) ;
assign n53 =  ( LB1D_p_cnt ) + ( 19'd1 )  ;
assign n54 =  ( 19'd316224 ) - ( 19'd1 )  ;
assign n55 =  ( LB1D_p_cnt ) == ( n54 )  ;
assign n56 =  ( n55 ) ? ( 19'd0 ) : ( n53 ) ;
assign n57 =  ( n37 ) ? ( n56 ) : ( LB1D_p_cnt ) ;
assign n58 =  ( n51 ) ? ( n53 ) : ( n57 ) ;
assign n59 =  ( n32 ) ? ( LB1D_p_cnt ) : ( n58 ) ;
assign n60 =  ( n25 ) ? ( LB1D_p_cnt ) : ( n59 ) ;
assign n61 =  ( n18 ) ? ( LB1D_p_cnt ) : ( n60 ) ;
assign n62 =  ( n9 ) ? ( LB1D_p_cnt ) : ( n61 ) ;
assign n63 =  ( n4 ) ? ( LB1D_p_cnt ) : ( n62 ) ;
assign n64 =  ( LB2D_proc_w ) < ( 64'd7 )  ;
assign n65 =  ( LB2D_proc_x ) < ( 9'd488 )  ;
assign n66 =  ( LB2D_proc_w ) + ( 64'd1 )  ;
assign n67 =  ( n65 ) ? ( LB2D_proc_w ) : ( n66 ) ;
assign n68 =  ( n64 ) ? ( n67 ) : ( 64'd0 ) ;
assign n69 =  ( n37 ) ? ( LB2D_proc_w ) : ( LB2D_proc_w ) ;
assign n70 =  ( n32 ) ? ( n68 ) : ( n69 ) ;
assign n71 =  ( n25 ) ? ( LB2D_proc_w ) : ( n70 ) ;
assign n72 =  ( n18 ) ? ( LB2D_proc_w ) : ( n71 ) ;
assign n73 =  ( n9 ) ? ( LB2D_proc_w ) : ( n72 ) ;
assign n74 =  ( n4 ) ? ( LB2D_proc_w ) : ( n73 ) ;
assign n75 =  ( LB2D_proc_x ) == ( 9'd488 )  ;
assign n76 =  ( n26 ) & ( n75 )  ;
assign n77 =  ( n76 ) & ( n31 )  ;
assign n78 =  ( LB2D_proc_x ) + ( 9'd1 )  ;
assign n79 =  ( n37 ) ? ( LB2D_proc_x ) : ( LB2D_proc_x ) ;
assign n80 =  ( n32 ) ? ( n78 ) : ( n79 ) ;
assign n81 =  ( n77 ) ? ( 9'd0 ) : ( n80 ) ;
assign n82 =  ( n25 ) ? ( LB2D_proc_x ) : ( n81 ) ;
assign n83 =  ( n18 ) ? ( LB2D_proc_x ) : ( n82 ) ;
assign n84 =  ( n9 ) ? ( LB2D_proc_x ) : ( n83 ) ;
assign n85 =  ( n4 ) ? ( LB2D_proc_x ) : ( n84 ) ;
assign n86 =  ( LB2D_proc_y ) < ( 10'd488 )  ;
assign n87 =  ( n86 ) ? ( LB2D_proc_y ) : ( 10'd488 ) ;
assign n88 =  ( n37 ) ? ( LB2D_proc_y ) : ( LB2D_proc_y ) ;
assign n89 =  ( n32 ) ? ( n87 ) : ( n88 ) ;
assign n90 =  ( n25 ) ? ( LB2D_proc_y ) : ( n89 ) ;
assign n91 =  ( n18 ) ? ( LB2D_proc_y ) : ( n90 ) ;
assign n92 =  ( n9 ) ? ( LB2D_proc_y ) : ( n91 ) ;
assign n93 =  ( n4 ) ? ( LB2D_proc_y ) : ( n92 ) ;
assign n94 =  ( slice_stream_full ) == ( 1'd1 )  ;
assign n95 =  ( n94 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n96 =  ( n37 ) ? ( LB2D_shift_0 ) : ( LB2D_shift_0 ) ;
assign n97 =  ( n32 ) ? ( LB2D_shift_0 ) : ( n96 ) ;
assign n98 =  ( n25 ) ? ( n95 ) : ( n97 ) ;
assign n99 =  ( n18 ) ? ( LB2D_shift_0 ) : ( n98 ) ;
assign n100 =  ( n9 ) ? ( LB2D_shift_0 ) : ( n99 ) ;
assign n101 =  ( n4 ) ? ( LB2D_shift_0 ) : ( n100 ) ;
assign n102 =  ( n37 ) ? ( LB2D_shift_1 ) : ( LB2D_shift_1 ) ;
assign n103 =  ( n32 ) ? ( LB2D_shift_1 ) : ( n102 ) ;
assign n104 =  ( n25 ) ? ( LB2D_shift_0 ) : ( n103 ) ;
assign n105 =  ( n18 ) ? ( LB2D_shift_1 ) : ( n104 ) ;
assign n106 =  ( n9 ) ? ( LB2D_shift_1 ) : ( n105 ) ;
assign n107 =  ( n4 ) ? ( LB2D_shift_1 ) : ( n106 ) ;
assign n108 =  ( n37 ) ? ( LB2D_shift_2 ) : ( LB2D_shift_2 ) ;
assign n109 =  ( n32 ) ? ( LB2D_shift_2 ) : ( n108 ) ;
assign n110 =  ( n25 ) ? ( LB2D_shift_1 ) : ( n109 ) ;
assign n111 =  ( n18 ) ? ( LB2D_shift_2 ) : ( n110 ) ;
assign n112 =  ( n9 ) ? ( LB2D_shift_2 ) : ( n111 ) ;
assign n113 =  ( n4 ) ? ( LB2D_shift_2 ) : ( n112 ) ;
assign n114 =  ( n37 ) ? ( LB2D_shift_3 ) : ( LB2D_shift_3 ) ;
assign n115 =  ( n32 ) ? ( LB2D_shift_3 ) : ( n114 ) ;
assign n116 =  ( n25 ) ? ( LB2D_shift_2 ) : ( n115 ) ;
assign n117 =  ( n18 ) ? ( LB2D_shift_3 ) : ( n116 ) ;
assign n118 =  ( n9 ) ? ( LB2D_shift_3 ) : ( n117 ) ;
assign n119 =  ( n4 ) ? ( LB2D_shift_3 ) : ( n118 ) ;
assign n120 =  ( n37 ) ? ( LB2D_shift_4 ) : ( LB2D_shift_4 ) ;
assign n121 =  ( n32 ) ? ( LB2D_shift_4 ) : ( n120 ) ;
assign n122 =  ( n25 ) ? ( LB2D_shift_3 ) : ( n121 ) ;
assign n123 =  ( n18 ) ? ( LB2D_shift_4 ) : ( n122 ) ;
assign n124 =  ( n9 ) ? ( LB2D_shift_4 ) : ( n123 ) ;
assign n125 =  ( n4 ) ? ( LB2D_shift_4 ) : ( n124 ) ;
assign n126 =  ( n37 ) ? ( LB2D_shift_5 ) : ( LB2D_shift_5 ) ;
assign n127 =  ( n32 ) ? ( LB2D_shift_5 ) : ( n126 ) ;
assign n128 =  ( n25 ) ? ( LB2D_shift_4 ) : ( n127 ) ;
assign n129 =  ( n18 ) ? ( LB2D_shift_5 ) : ( n128 ) ;
assign n130 =  ( n9 ) ? ( LB2D_shift_5 ) : ( n129 ) ;
assign n131 =  ( n4 ) ? ( LB2D_shift_5 ) : ( n130 ) ;
assign n132 =  ( n37 ) ? ( LB2D_shift_6 ) : ( LB2D_shift_6 ) ;
assign n133 =  ( n32 ) ? ( LB2D_shift_6 ) : ( n132 ) ;
assign n134 =  ( n25 ) ? ( LB2D_shift_5 ) : ( n133 ) ;
assign n135 =  ( n18 ) ? ( LB2D_shift_6 ) : ( n134 ) ;
assign n136 =  ( n9 ) ? ( LB2D_shift_6 ) : ( n135 ) ;
assign n137 =  ( n4 ) ? ( LB2D_shift_6 ) : ( n136 ) ;
assign n138 =  ( n37 ) ? ( LB2D_shift_7 ) : ( LB2D_shift_7 ) ;
assign n139 =  ( n32 ) ? ( LB2D_shift_7 ) : ( n138 ) ;
assign n140 =  ( n25 ) ? ( LB2D_shift_6 ) : ( n139 ) ;
assign n141 =  ( n18 ) ? ( LB2D_shift_7 ) : ( n140 ) ;
assign n142 =  ( n9 ) ? ( LB2D_shift_7 ) : ( n141 ) ;
assign n143 =  ( n4 ) ? ( LB2D_shift_7 ) : ( n142 ) ;
assign n144 =  ( LB2D_shift_x ) + ( 9'd1 )  ;
assign n145 =  ( n37 ) ? ( LB2D_shift_x ) : ( LB2D_shift_x ) ;
assign n146 =  ( n32 ) ? ( LB2D_shift_x ) : ( n145 ) ;
assign n147 =  ( n25 ) ? ( n144 ) : ( n146 ) ;
assign n148 =  ( n18 ) ? ( LB2D_shift_x ) : ( n147 ) ;
assign n149 =  ( n9 ) ? ( LB2D_shift_x ) : ( n148 ) ;
assign n150 =  ( n4 ) ? ( LB2D_shift_x ) : ( n149 ) ;
assign n151 =  ( LB2D_shift_y ) < ( 10'd480 )  ;
assign n152 =  ( LB2D_shift_x ) < ( 9'd488 )  ;
assign n153 =  ( LB2D_shift_y ) + ( 10'd1 )  ;
assign n154 =  ( n152 ) ? ( LB2D_shift_y ) : ( n153 ) ;
assign n155 =  ( n151 ) ? ( n154 ) : ( 10'd480 ) ;
assign n156 =  ( n37 ) ? ( LB2D_shift_y ) : ( LB2D_shift_y ) ;
assign n157 =  ( n32 ) ? ( LB2D_shift_y ) : ( n156 ) ;
assign n158 =  ( n25 ) ? ( n155 ) : ( n157 ) ;
assign n159 =  ( n18 ) ? ( LB2D_shift_y ) : ( n158 ) ;
assign n160 =  ( n9 ) ? ( LB2D_shift_y ) : ( n159 ) ;
assign n161 =  ( n4 ) ? ( LB2D_shift_y ) : ( n160 ) ;
assign n162 =  ( stencil_stream_full ) == ( 1'd1 )  ;
assign n163 =  ( n162 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_0 ) ;
assign n164 = gb_fun(n163) ;
assign n165 =  ( n37 ) ? ( arg_0_TDATA ) : ( arg_0_TDATA ) ;
assign n166 =  ( n32 ) ? ( arg_0_TDATA ) : ( n165 ) ;
assign n167 =  ( n25 ) ? ( arg_0_TDATA ) : ( n166 ) ;
assign n168 =  ( n18 ) ? ( n164 ) : ( n167 ) ;
assign n169 =  ( n9 ) ? ( arg_0_TDATA ) : ( n168 ) ;
assign n170 =  ( n4 ) ? ( arg_0_TDATA ) : ( n169 ) ;
assign n171 =  ( gb_pp_it_8 ) == ( 1'd1 )  ;
assign n172 =  ( n171 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n173 =  ( n37 ) ? ( arg_0_TVALID ) : ( arg_0_TVALID ) ;
assign n174 =  ( n32 ) ? ( arg_0_TVALID ) : ( n173 ) ;
assign n175 =  ( n25 ) ? ( arg_0_TVALID ) : ( n174 ) ;
assign n176 =  ( n18 ) ? ( n172 ) : ( n175 ) ;
assign n177 =  ( n9 ) ? ( arg_0_TVALID ) : ( n176 ) ;
assign n178 =  ( n4 ) ? ( 1'd0 ) : ( n177 ) ;
assign n179 =  ( n37 ) ? ( 1'd1 ) : ( arg_1_TREADY ) ;
assign n180 =  ( n51 ) ? ( 1'd1 ) : ( n179 ) ;
assign n181 =  ( n32 ) ? ( arg_1_TREADY ) : ( n180 ) ;
assign n182 =  ( n25 ) ? ( arg_1_TREADY ) : ( n181 ) ;
assign n183 =  ( n18 ) ? ( arg_1_TREADY ) : ( n182 ) ;
assign n184 =  ( n9 ) ? ( 1'd0 ) : ( n183 ) ;
assign n185 =  ( n4 ) ? ( 1'd0 ) : ( n184 ) ;
assign n186 =  ( gb_p_cnt ) + ( 19'd1 )  ;
assign n187 =  ( n186 ) == ( 19'd307200 )  ;
assign n188 =  ( n187 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n189 =  ( n37 ) ? ( gb_exit_it_1 ) : ( gb_exit_it_1 ) ;
assign n190 =  ( n32 ) ? ( gb_exit_it_1 ) : ( n189 ) ;
assign n191 =  ( n25 ) ? ( gb_exit_it_1 ) : ( n190 ) ;
assign n192 =  ( n18 ) ? ( n188 ) : ( n191 ) ;
assign n193 =  ( n9 ) ? ( gb_exit_it_1 ) : ( n192 ) ;
assign n194 =  ( n4 ) ? ( gb_exit_it_1 ) : ( n193 ) ;
assign n195 =  ( n37 ) ? ( gb_exit_it_2 ) : ( gb_exit_it_2 ) ;
assign n196 =  ( n32 ) ? ( gb_exit_it_2 ) : ( n195 ) ;
assign n197 =  ( n25 ) ? ( gb_exit_it_2 ) : ( n196 ) ;
assign n198 =  ( n18 ) ? ( gb_exit_it_1 ) : ( n197 ) ;
assign n199 =  ( n9 ) ? ( gb_exit_it_2 ) : ( n198 ) ;
assign n200 =  ( n4 ) ? ( gb_exit_it_2 ) : ( n199 ) ;
assign n201 =  ( n37 ) ? ( gb_exit_it_3 ) : ( gb_exit_it_3 ) ;
assign n202 =  ( n32 ) ? ( gb_exit_it_3 ) : ( n201 ) ;
assign n203 =  ( n25 ) ? ( gb_exit_it_3 ) : ( n202 ) ;
assign n204 =  ( n18 ) ? ( gb_exit_it_2 ) : ( n203 ) ;
assign n205 =  ( n9 ) ? ( gb_exit_it_3 ) : ( n204 ) ;
assign n206 =  ( n4 ) ? ( gb_exit_it_3 ) : ( n205 ) ;
assign n207 =  ( n37 ) ? ( gb_exit_it_4 ) : ( gb_exit_it_4 ) ;
assign n208 =  ( n32 ) ? ( gb_exit_it_4 ) : ( n207 ) ;
assign n209 =  ( n25 ) ? ( gb_exit_it_4 ) : ( n208 ) ;
assign n210 =  ( n18 ) ? ( gb_exit_it_3 ) : ( n209 ) ;
assign n211 =  ( n9 ) ? ( gb_exit_it_4 ) : ( n210 ) ;
assign n212 =  ( n4 ) ? ( gb_exit_it_4 ) : ( n211 ) ;
assign n213 =  ( n37 ) ? ( gb_exit_it_5 ) : ( gb_exit_it_5 ) ;
assign n214 =  ( n32 ) ? ( gb_exit_it_5 ) : ( n213 ) ;
assign n215 =  ( n25 ) ? ( gb_exit_it_5 ) : ( n214 ) ;
assign n216 =  ( n18 ) ? ( gb_exit_it_4 ) : ( n215 ) ;
assign n217 =  ( n9 ) ? ( gb_exit_it_5 ) : ( n216 ) ;
assign n218 =  ( n4 ) ? ( gb_exit_it_5 ) : ( n217 ) ;
assign n219 =  ( n37 ) ? ( gb_exit_it_6 ) : ( gb_exit_it_6 ) ;
assign n220 =  ( n32 ) ? ( gb_exit_it_6 ) : ( n219 ) ;
assign n221 =  ( n25 ) ? ( gb_exit_it_6 ) : ( n220 ) ;
assign n222 =  ( n18 ) ? ( gb_exit_it_5 ) : ( n221 ) ;
assign n223 =  ( n9 ) ? ( gb_exit_it_6 ) : ( n222 ) ;
assign n224 =  ( n4 ) ? ( gb_exit_it_6 ) : ( n223 ) ;
assign n225 =  ( n37 ) ? ( gb_exit_it_7 ) : ( gb_exit_it_7 ) ;
assign n226 =  ( n32 ) ? ( gb_exit_it_7 ) : ( n225 ) ;
assign n227 =  ( n25 ) ? ( gb_exit_it_7 ) : ( n226 ) ;
assign n228 =  ( n18 ) ? ( gb_exit_it_6 ) : ( n227 ) ;
assign n229 =  ( n9 ) ? ( gb_exit_it_7 ) : ( n228 ) ;
assign n230 =  ( n4 ) ? ( gb_exit_it_7 ) : ( n229 ) ;
assign n231 =  ( n37 ) ? ( gb_exit_it_8 ) : ( gb_exit_it_8 ) ;
assign n232 =  ( n32 ) ? ( gb_exit_it_8 ) : ( n231 ) ;
assign n233 =  ( n25 ) ? ( gb_exit_it_8 ) : ( n232 ) ;
assign n234 =  ( n18 ) ? ( gb_exit_it_7 ) : ( n233 ) ;
assign n235 =  ( n9 ) ? ( gb_exit_it_8 ) : ( n234 ) ;
assign n236 =  ( n4 ) ? ( gb_exit_it_8 ) : ( n235 ) ;
assign n237 =  ( gb_p_cnt ) < ( 19'd307200 )  ;
assign n238 =  ( n237 ) ? ( n186 ) : ( 19'd307200 ) ;
assign n239 =  ( n37 ) ? ( gb_p_cnt ) : ( gb_p_cnt ) ;
assign n240 =  ( n32 ) ? ( gb_p_cnt ) : ( n239 ) ;
assign n241 =  ( n25 ) ? ( gb_p_cnt ) : ( n240 ) ;
assign n242 =  ( n18 ) ? ( n238 ) : ( n241 ) ;
assign n243 =  ( n9 ) ? ( gb_p_cnt ) : ( n242 ) ;
assign n244 =  ( n4 ) ? ( gb_p_cnt ) : ( n243 ) ;
assign n245 =  ( n37 ) ? ( gb_pp_it_1 ) : ( gb_pp_it_1 ) ;
assign n246 =  ( n32 ) ? ( gb_pp_it_1 ) : ( n245 ) ;
assign n247 =  ( n25 ) ? ( gb_pp_it_1 ) : ( n246 ) ;
assign n248 =  ( n18 ) ? ( 1'd1 ) : ( n247 ) ;
assign n249 =  ( n9 ) ? ( gb_pp_it_1 ) : ( n248 ) ;
assign n250 =  ( n4 ) ? ( gb_pp_it_1 ) : ( n249 ) ;
assign n251 =  ( n37 ) ? ( gb_pp_it_2 ) : ( gb_pp_it_2 ) ;
assign n252 =  ( n32 ) ? ( gb_pp_it_2 ) : ( n251 ) ;
assign n253 =  ( n25 ) ? ( gb_pp_it_2 ) : ( n252 ) ;
assign n254 =  ( n18 ) ? ( gb_pp_it_1 ) : ( n253 ) ;
assign n255 =  ( n9 ) ? ( gb_pp_it_2 ) : ( n254 ) ;
assign n256 =  ( n4 ) ? ( gb_pp_it_2 ) : ( n255 ) ;
assign n257 =  ( n37 ) ? ( gb_pp_it_3 ) : ( gb_pp_it_3 ) ;
assign n258 =  ( n32 ) ? ( gb_pp_it_3 ) : ( n257 ) ;
assign n259 =  ( n25 ) ? ( gb_pp_it_3 ) : ( n258 ) ;
assign n260 =  ( n18 ) ? ( gb_pp_it_2 ) : ( n259 ) ;
assign n261 =  ( n9 ) ? ( gb_pp_it_3 ) : ( n260 ) ;
assign n262 =  ( n4 ) ? ( gb_pp_it_3 ) : ( n261 ) ;
assign n263 =  ( n37 ) ? ( gb_pp_it_4 ) : ( gb_pp_it_4 ) ;
assign n264 =  ( n32 ) ? ( gb_pp_it_4 ) : ( n263 ) ;
assign n265 =  ( n25 ) ? ( gb_pp_it_4 ) : ( n264 ) ;
assign n266 =  ( n18 ) ? ( gb_pp_it_3 ) : ( n265 ) ;
assign n267 =  ( n9 ) ? ( gb_pp_it_4 ) : ( n266 ) ;
assign n268 =  ( n4 ) ? ( gb_pp_it_4 ) : ( n267 ) ;
assign n269 =  ( n37 ) ? ( gb_pp_it_5 ) : ( gb_pp_it_5 ) ;
assign n270 =  ( n32 ) ? ( gb_pp_it_5 ) : ( n269 ) ;
assign n271 =  ( n25 ) ? ( gb_pp_it_5 ) : ( n270 ) ;
assign n272 =  ( n18 ) ? ( gb_pp_it_4 ) : ( n271 ) ;
assign n273 =  ( n9 ) ? ( gb_pp_it_5 ) : ( n272 ) ;
assign n274 =  ( n4 ) ? ( gb_pp_it_5 ) : ( n273 ) ;
assign n275 =  ( n37 ) ? ( gb_pp_it_6 ) : ( gb_pp_it_6 ) ;
assign n276 =  ( n32 ) ? ( gb_pp_it_6 ) : ( n275 ) ;
assign n277 =  ( n25 ) ? ( gb_pp_it_6 ) : ( n276 ) ;
assign n278 =  ( n18 ) ? ( gb_pp_it_5 ) : ( n277 ) ;
assign n279 =  ( n9 ) ? ( gb_pp_it_6 ) : ( n278 ) ;
assign n280 =  ( n4 ) ? ( gb_pp_it_6 ) : ( n279 ) ;
assign n281 =  ( n37 ) ? ( gb_pp_it_7 ) : ( gb_pp_it_7 ) ;
assign n282 =  ( n32 ) ? ( gb_pp_it_7 ) : ( n281 ) ;
assign n283 =  ( n25 ) ? ( gb_pp_it_7 ) : ( n282 ) ;
assign n284 =  ( n18 ) ? ( gb_pp_it_6 ) : ( n283 ) ;
assign n285 =  ( n9 ) ? ( gb_pp_it_7 ) : ( n284 ) ;
assign n286 =  ( n4 ) ? ( gb_pp_it_7 ) : ( n285 ) ;
assign n287 =  ( n37 ) ? ( gb_pp_it_8 ) : ( gb_pp_it_8 ) ;
assign n288 =  ( n32 ) ? ( gb_pp_it_8 ) : ( n287 ) ;
assign n289 =  ( n25 ) ? ( gb_pp_it_8 ) : ( n288 ) ;
assign n290 =  ( n18 ) ? ( gb_pp_it_7 ) : ( n289 ) ;
assign n291 =  ( n9 ) ? ( gb_pp_it_8 ) : ( n290 ) ;
assign n292 =  ( n4 ) ? ( gb_pp_it_8 ) : ( n291 ) ;
assign n293 =  ( n37 ) ? ( gb_pp_it_9 ) : ( gb_pp_it_9 ) ;
assign n294 =  ( n32 ) ? ( gb_pp_it_9 ) : ( n293 ) ;
assign n295 =  ( n25 ) ? ( gb_pp_it_9 ) : ( n294 ) ;
assign n296 =  ( n18 ) ? ( gb_pp_it_8 ) : ( n295 ) ;
assign n297 =  ( n9 ) ? ( gb_pp_it_9 ) : ( n296 ) ;
assign n298 =  ( n4 ) ? ( gb_pp_it_9 ) : ( n297 ) ;
assign n299 =  ( n37 ) ? ( LB1D_buff ) : ( in_stream_buff_0 ) ;
assign n300 =  ( n32 ) ? ( in_stream_buff_0 ) : ( n299 ) ;
assign n301 =  ( n25 ) ? ( in_stream_buff_0 ) : ( n300 ) ;
assign n302 =  ( n18 ) ? ( in_stream_buff_0 ) : ( n301 ) ;
assign n303 =  ( n9 ) ? ( in_stream_buff_0 ) : ( n302 ) ;
assign n304 =  ( n4 ) ? ( in_stream_buff_0 ) : ( n303 ) ;
assign n305 =  ( n37 ) ? ( in_stream_buff_0 ) : ( in_stream_buff_1 ) ;
assign n306 =  ( n32 ) ? ( in_stream_buff_1 ) : ( n305 ) ;
assign n307 =  ( n25 ) ? ( in_stream_buff_1 ) : ( n306 ) ;
assign n308 =  ( n18 ) ? ( in_stream_buff_1 ) : ( n307 ) ;
assign n309 =  ( n9 ) ? ( in_stream_buff_1 ) : ( n308 ) ;
assign n310 =  ( n4 ) ? ( in_stream_buff_1 ) : ( n309 ) ;
assign n311 =  ( in_stream_full ) == ( 1'd1 )  ;
assign n312 =  ( n311 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n313 =  ( n37 ) ? ( 1'd0 ) : ( in_stream_empty ) ;
assign n314 =  ( n32 ) ? ( n312 ) : ( n313 ) ;
assign n315 =  ( n25 ) ? ( in_stream_empty ) : ( n314 ) ;
assign n316 =  ( n18 ) ? ( in_stream_empty ) : ( n315 ) ;
assign n317 =  ( n9 ) ? ( in_stream_empty ) : ( n316 ) ;
assign n318 =  ( n4 ) ? ( in_stream_empty ) : ( n317 ) ;
assign n319 =  ( in_stream_empty ) == ( 1'd1 )  ;
assign n320 =  ( n319 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n321 =  ( n37 ) ? ( n320 ) : ( in_stream_full ) ;
assign n322 =  ( n32 ) ? ( 1'd0 ) : ( n321 ) ;
assign n323 =  ( n25 ) ? ( in_stream_full ) : ( n322 ) ;
assign n324 =  ( n18 ) ? ( in_stream_full ) : ( n323 ) ;
assign n325 =  ( n9 ) ? ( in_stream_full ) : ( n324 ) ;
assign n326 =  ( n4 ) ? ( in_stream_full ) : ( n325 ) ;
assign n327 =  ( n311 ) ? ( in_stream_buff_1 ) : ( in_stream_buff_0 ) ;
assign n328 =  ( LB2D_proc_w ) == ( 64'd0 )  ;
assign n329 =  (  LB2D_proc_7 [ LB2D_proc_x ] )  ;
assign n330 =  ( LB2D_proc_w ) == ( 64'd1 )  ;
assign n331 =  (  LB2D_proc_0 [ LB2D_proc_x ] )  ;
assign n332 =  ( LB2D_proc_w ) == ( 64'd2 )  ;
assign n333 =  (  LB2D_proc_1 [ LB2D_proc_x ] )  ;
assign n334 =  ( LB2D_proc_w ) == ( 64'd3 )  ;
assign n335 =  (  LB2D_proc_2 [ LB2D_proc_x ] )  ;
assign n336 =  ( LB2D_proc_w ) == ( 64'd4 )  ;
assign n337 =  (  LB2D_proc_3 [ LB2D_proc_x ] )  ;
assign n338 =  ( LB2D_proc_w ) == ( 64'd5 )  ;
assign n339 =  (  LB2D_proc_4 [ LB2D_proc_x ] )  ;
assign n340 =  ( LB2D_proc_w ) == ( 64'd6 )  ;
assign n341 =  (  LB2D_proc_5 [ LB2D_proc_x ] )  ;
assign n342 =  (  LB2D_proc_6 [ LB2D_proc_x ] )  ;
assign n343 =  ( n340 ) ? ( n341 ) : ( n342 ) ;
assign n344 =  ( n338 ) ? ( n339 ) : ( n343 ) ;
assign n345 =  ( n336 ) ? ( n337 ) : ( n344 ) ;
assign n346 =  ( n334 ) ? ( n335 ) : ( n345 ) ;
assign n347 =  ( n332 ) ? ( n333 ) : ( n346 ) ;
assign n348 =  ( n330 ) ? ( n331 ) : ( n347 ) ;
assign n349 =  ( n328 ) ? ( n329 ) : ( n348 ) ;
assign n350 =  ( n340 ) ? ( n339 ) : ( n341 ) ;
assign n351 =  ( n338 ) ? ( n337 ) : ( n350 ) ;
assign n352 =  ( n336 ) ? ( n335 ) : ( n351 ) ;
assign n353 =  ( n334 ) ? ( n333 ) : ( n352 ) ;
assign n354 =  ( n332 ) ? ( n331 ) : ( n353 ) ;
assign n355 =  ( n330 ) ? ( n329 ) : ( n354 ) ;
assign n356 =  ( n328 ) ? ( n342 ) : ( n355 ) ;
assign n357 =  ( n340 ) ? ( n337 ) : ( n339 ) ;
assign n358 =  ( n338 ) ? ( n335 ) : ( n357 ) ;
assign n359 =  ( n336 ) ? ( n333 ) : ( n358 ) ;
assign n360 =  ( n334 ) ? ( n331 ) : ( n359 ) ;
assign n361 =  ( n332 ) ? ( n329 ) : ( n360 ) ;
assign n362 =  ( n330 ) ? ( n342 ) : ( n361 ) ;
assign n363 =  ( n328 ) ? ( n341 ) : ( n362 ) ;
assign n364 =  ( n340 ) ? ( n335 ) : ( n337 ) ;
assign n365 =  ( n338 ) ? ( n333 ) : ( n364 ) ;
assign n366 =  ( n336 ) ? ( n331 ) : ( n365 ) ;
assign n367 =  ( n334 ) ? ( n329 ) : ( n366 ) ;
assign n368 =  ( n332 ) ? ( n342 ) : ( n367 ) ;
assign n369 =  ( n330 ) ? ( n341 ) : ( n368 ) ;
assign n370 =  ( n328 ) ? ( n339 ) : ( n369 ) ;
assign n371 =  ( n340 ) ? ( n333 ) : ( n335 ) ;
assign n372 =  ( n338 ) ? ( n331 ) : ( n371 ) ;
assign n373 =  ( n336 ) ? ( n329 ) : ( n372 ) ;
assign n374 =  ( n334 ) ? ( n342 ) : ( n373 ) ;
assign n375 =  ( n332 ) ? ( n341 ) : ( n374 ) ;
assign n376 =  ( n330 ) ? ( n339 ) : ( n375 ) ;
assign n377 =  ( n328 ) ? ( n337 ) : ( n376 ) ;
assign n378 =  ( n340 ) ? ( n331 ) : ( n333 ) ;
assign n379 =  ( n338 ) ? ( n329 ) : ( n378 ) ;
assign n380 =  ( n336 ) ? ( n342 ) : ( n379 ) ;
assign n381 =  ( n334 ) ? ( n341 ) : ( n380 ) ;
assign n382 =  ( n332 ) ? ( n339 ) : ( n381 ) ;
assign n383 =  ( n330 ) ? ( n337 ) : ( n382 ) ;
assign n384 =  ( n328 ) ? ( n335 ) : ( n383 ) ;
assign n385 =  ( n340 ) ? ( n329 ) : ( n331 ) ;
assign n386 =  ( n338 ) ? ( n342 ) : ( n385 ) ;
assign n387 =  ( n336 ) ? ( n341 ) : ( n386 ) ;
assign n388 =  ( n334 ) ? ( n339 ) : ( n387 ) ;
assign n389 =  ( n332 ) ? ( n337 ) : ( n388 ) ;
assign n390 =  ( n330 ) ? ( n335 ) : ( n389 ) ;
assign n391 =  ( n328 ) ? ( n333 ) : ( n390 ) ;
assign n392 =  ( n340 ) ? ( n342 ) : ( n329 ) ;
assign n393 =  ( n338 ) ? ( n341 ) : ( n392 ) ;
assign n394 =  ( n336 ) ? ( n339 ) : ( n393 ) ;
assign n395 =  ( n334 ) ? ( n337 ) : ( n394 ) ;
assign n396 =  ( n332 ) ? ( n335 ) : ( n395 ) ;
assign n397 =  ( n330 ) ? ( n333 ) : ( n396 ) ;
assign n398 =  ( n328 ) ? ( n331 ) : ( n397 ) ;
assign n399 =  { ( n391 ) , ( n398 ) }  ;
assign n400 =  { ( n384 ) , ( n399 ) }  ;
assign n401 =  { ( n377 ) , ( n400 ) }  ;
assign n402 =  { ( n370 ) , ( n401 ) }  ;
assign n403 =  { ( n363 ) , ( n402 ) }  ;
assign n404 =  { ( n356 ) , ( n403 ) }  ;
assign n405 =  { ( n349 ) , ( n404 ) }  ;
assign n406 =  { ( n327 ) , ( n405 ) }  ;
assign n407 =  ( n30 ) ? ( slice_stream_buff_0 ) : ( n406 ) ;
assign n408 =  ( n37 ) ? ( slice_stream_buff_0 ) : ( slice_stream_buff_0 ) ;
assign n409 =  ( n32 ) ? ( n407 ) : ( n408 ) ;
assign n410 =  ( n25 ) ? ( slice_stream_buff_0 ) : ( n409 ) ;
assign n411 =  ( n18 ) ? ( slice_stream_buff_0 ) : ( n410 ) ;
assign n412 =  ( n9 ) ? ( slice_stream_buff_0 ) : ( n411 ) ;
assign n413 =  ( n4 ) ? ( slice_stream_buff_0 ) : ( n412 ) ;
assign n414 =  ( n30 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n415 =  ( n37 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_1 ) ;
assign n416 =  ( n32 ) ? ( n414 ) : ( n415 ) ;
assign n417 =  ( n25 ) ? ( slice_stream_buff_1 ) : ( n416 ) ;
assign n418 =  ( n18 ) ? ( slice_stream_buff_1 ) : ( n417 ) ;
assign n419 =  ( n9 ) ? ( slice_stream_buff_1 ) : ( n418 ) ;
assign n420 =  ( n4 ) ? ( slice_stream_buff_1 ) : ( n419 ) ;
assign n421 =  ( n94 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n422 =  ( n30 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n423 =  ( n37 ) ? ( slice_stream_empty ) : ( slice_stream_empty ) ;
assign n424 =  ( n32 ) ? ( n422 ) : ( n423 ) ;
assign n425 =  ( n25 ) ? ( n421 ) : ( n424 ) ;
assign n426 =  ( n18 ) ? ( slice_stream_empty ) : ( n425 ) ;
assign n427 =  ( n9 ) ? ( slice_stream_empty ) : ( n426 ) ;
assign n428 =  ( n4 ) ? ( slice_stream_empty ) : ( n427 ) ;
assign n429 =  ( slice_stream_empty ) == ( 1'd1 )  ;
assign n430 =  ( n429 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n431 =  ( n30 ) ? ( 1'd0 ) : ( n430 ) ;
assign n432 =  ( n37 ) ? ( slice_stream_full ) : ( slice_stream_full ) ;
assign n433 =  ( n32 ) ? ( n431 ) : ( n432 ) ;
assign n434 =  ( n25 ) ? ( 1'd0 ) : ( n433 ) ;
assign n435 =  ( n18 ) ? ( slice_stream_full ) : ( n434 ) ;
assign n436 =  ( n9 ) ? ( slice_stream_full ) : ( n435 ) ;
assign n437 =  ( n4 ) ? ( slice_stream_full ) : ( n436 ) ;
assign n438 =  ( LB2D_shift_x ) >= ( 9'd8 )  ;
assign n439 = n95[71:64] ;
assign n440 = LB2D_shift_0[71:64] ;
assign n441 = LB2D_shift_1[71:64] ;
assign n442 = LB2D_shift_2[71:64] ;
assign n443 = LB2D_shift_3[71:64] ;
assign n444 = LB2D_shift_4[71:64] ;
assign n445 = LB2D_shift_5[71:64] ;
assign n446 = LB2D_shift_6[71:64] ;
assign n447 = LB2D_shift_7[71:64] ;
assign n448 =  { ( n446 ) , ( n447 ) }  ;
assign n449 =  { ( n445 ) , ( n448 ) }  ;
assign n450 =  { ( n444 ) , ( n449 ) }  ;
assign n451 =  { ( n443 ) , ( n450 ) }  ;
assign n452 =  { ( n442 ) , ( n451 ) }  ;
assign n453 =  { ( n441 ) , ( n452 ) }  ;
assign n454 =  { ( n440 ) , ( n453 ) }  ;
assign n455 =  { ( n439 ) , ( n454 ) }  ;
assign n456 = n95[63:56] ;
assign n457 = LB2D_shift_0[63:56] ;
assign n458 = LB2D_shift_1[63:56] ;
assign n459 = LB2D_shift_2[63:56] ;
assign n460 = LB2D_shift_3[63:56] ;
assign n461 = LB2D_shift_4[63:56] ;
assign n462 = LB2D_shift_5[63:56] ;
assign n463 = LB2D_shift_6[63:56] ;
assign n464 = LB2D_shift_7[63:56] ;
assign n465 =  { ( n463 ) , ( n464 ) }  ;
assign n466 =  { ( n462 ) , ( n465 ) }  ;
assign n467 =  { ( n461 ) , ( n466 ) }  ;
assign n468 =  { ( n460 ) , ( n467 ) }  ;
assign n469 =  { ( n459 ) , ( n468 ) }  ;
assign n470 =  { ( n458 ) , ( n469 ) }  ;
assign n471 =  { ( n457 ) , ( n470 ) }  ;
assign n472 =  { ( n456 ) , ( n471 ) }  ;
assign n473 = n95[55:48] ;
assign n474 = LB2D_shift_0[55:48] ;
assign n475 = LB2D_shift_1[55:48] ;
assign n476 = LB2D_shift_2[55:48] ;
assign n477 = LB2D_shift_3[55:48] ;
assign n478 = LB2D_shift_4[55:48] ;
assign n479 = LB2D_shift_5[55:48] ;
assign n480 = LB2D_shift_6[55:48] ;
assign n481 = LB2D_shift_7[55:48] ;
assign n482 =  { ( n480 ) , ( n481 ) }  ;
assign n483 =  { ( n479 ) , ( n482 ) }  ;
assign n484 =  { ( n478 ) , ( n483 ) }  ;
assign n485 =  { ( n477 ) , ( n484 ) }  ;
assign n486 =  { ( n476 ) , ( n485 ) }  ;
assign n487 =  { ( n475 ) , ( n486 ) }  ;
assign n488 =  { ( n474 ) , ( n487 ) }  ;
assign n489 =  { ( n473 ) , ( n488 ) }  ;
assign n490 = n95[47:40] ;
assign n491 = LB2D_shift_0[47:40] ;
assign n492 = LB2D_shift_1[47:40] ;
assign n493 = LB2D_shift_2[47:40] ;
assign n494 = LB2D_shift_3[47:40] ;
assign n495 = LB2D_shift_4[47:40] ;
assign n496 = LB2D_shift_5[47:40] ;
assign n497 = LB2D_shift_6[47:40] ;
assign n498 = LB2D_shift_7[47:40] ;
assign n499 =  { ( n497 ) , ( n498 ) }  ;
assign n500 =  { ( n496 ) , ( n499 ) }  ;
assign n501 =  { ( n495 ) , ( n500 ) }  ;
assign n502 =  { ( n494 ) , ( n501 ) }  ;
assign n503 =  { ( n493 ) , ( n502 ) }  ;
assign n504 =  { ( n492 ) , ( n503 ) }  ;
assign n505 =  { ( n491 ) , ( n504 ) }  ;
assign n506 =  { ( n490 ) , ( n505 ) }  ;
assign n507 = n95[39:32] ;
assign n508 = LB2D_shift_0[39:32] ;
assign n509 = LB2D_shift_1[39:32] ;
assign n510 = LB2D_shift_2[39:32] ;
assign n511 = LB2D_shift_3[39:32] ;
assign n512 = LB2D_shift_4[39:32] ;
assign n513 = LB2D_shift_5[39:32] ;
assign n514 = LB2D_shift_6[39:32] ;
assign n515 = LB2D_shift_7[39:32] ;
assign n516 =  { ( n514 ) , ( n515 ) }  ;
assign n517 =  { ( n513 ) , ( n516 ) }  ;
assign n518 =  { ( n512 ) , ( n517 ) }  ;
assign n519 =  { ( n511 ) , ( n518 ) }  ;
assign n520 =  { ( n510 ) , ( n519 ) }  ;
assign n521 =  { ( n509 ) , ( n520 ) }  ;
assign n522 =  { ( n508 ) , ( n521 ) }  ;
assign n523 =  { ( n507 ) , ( n522 ) }  ;
assign n524 = n95[31:24] ;
assign n525 = LB2D_shift_0[31:24] ;
assign n526 = LB2D_shift_1[31:24] ;
assign n527 = LB2D_shift_2[31:24] ;
assign n528 = LB2D_shift_3[31:24] ;
assign n529 = LB2D_shift_4[31:24] ;
assign n530 = LB2D_shift_5[31:24] ;
assign n531 = LB2D_shift_6[31:24] ;
assign n532 = LB2D_shift_7[31:24] ;
assign n533 =  { ( n531 ) , ( n532 ) }  ;
assign n534 =  { ( n530 ) , ( n533 ) }  ;
assign n535 =  { ( n529 ) , ( n534 ) }  ;
assign n536 =  { ( n528 ) , ( n535 ) }  ;
assign n537 =  { ( n527 ) , ( n536 ) }  ;
assign n538 =  { ( n526 ) , ( n537 ) }  ;
assign n539 =  { ( n525 ) , ( n538 ) }  ;
assign n540 =  { ( n524 ) , ( n539 ) }  ;
assign n541 = n95[23:16] ;
assign n542 = LB2D_shift_0[23:16] ;
assign n543 = LB2D_shift_1[23:16] ;
assign n544 = LB2D_shift_2[23:16] ;
assign n545 = LB2D_shift_3[23:16] ;
assign n546 = LB2D_shift_4[23:16] ;
assign n547 = LB2D_shift_5[23:16] ;
assign n548 = LB2D_shift_6[23:16] ;
assign n549 = LB2D_shift_7[23:16] ;
assign n550 =  { ( n548 ) , ( n549 ) }  ;
assign n551 =  { ( n547 ) , ( n550 ) }  ;
assign n552 =  { ( n546 ) , ( n551 ) }  ;
assign n553 =  { ( n545 ) , ( n552 ) }  ;
assign n554 =  { ( n544 ) , ( n553 ) }  ;
assign n555 =  { ( n543 ) , ( n554 ) }  ;
assign n556 =  { ( n542 ) , ( n555 ) }  ;
assign n557 =  { ( n541 ) , ( n556 ) }  ;
assign n558 = n95[15:8] ;
assign n559 = LB2D_shift_0[15:8] ;
assign n560 = LB2D_shift_1[15:8] ;
assign n561 = LB2D_shift_2[15:8] ;
assign n562 = LB2D_shift_3[15:8] ;
assign n563 = LB2D_shift_4[15:8] ;
assign n564 = LB2D_shift_5[15:8] ;
assign n565 = LB2D_shift_6[15:8] ;
assign n566 = LB2D_shift_7[15:8] ;
assign n567 =  { ( n565 ) , ( n566 ) }  ;
assign n568 =  { ( n564 ) , ( n567 ) }  ;
assign n569 =  { ( n563 ) , ( n568 ) }  ;
assign n570 =  { ( n562 ) , ( n569 ) }  ;
assign n571 =  { ( n561 ) , ( n570 ) }  ;
assign n572 =  { ( n560 ) , ( n571 ) }  ;
assign n573 =  { ( n559 ) , ( n572 ) }  ;
assign n574 =  { ( n558 ) , ( n573 ) }  ;
assign n575 = n95[7:0] ;
assign n576 = LB2D_shift_0[7:0] ;
assign n577 = LB2D_shift_1[7:0] ;
assign n578 = LB2D_shift_2[7:0] ;
assign n579 = LB2D_shift_3[7:0] ;
assign n580 = LB2D_shift_4[7:0] ;
assign n581 = LB2D_shift_5[7:0] ;
assign n582 = LB2D_shift_6[7:0] ;
assign n583 = LB2D_shift_7[7:0] ;
assign n584 =  { ( n582 ) , ( n583 ) }  ;
assign n585 =  { ( n581 ) , ( n584 ) }  ;
assign n586 =  { ( n580 ) , ( n585 ) }  ;
assign n587 =  { ( n579 ) , ( n586 ) }  ;
assign n588 =  { ( n578 ) , ( n587 ) }  ;
assign n589 =  { ( n577 ) , ( n588 ) }  ;
assign n590 =  { ( n576 ) , ( n589 ) }  ;
assign n591 =  { ( n575 ) , ( n590 ) }  ;
assign n592 =  { ( n574 ) , ( n591 ) }  ;
assign n593 =  { ( n557 ) , ( n592 ) }  ;
assign n594 =  { ( n540 ) , ( n593 ) }  ;
assign n595 =  { ( n523 ) , ( n594 ) }  ;
assign n596 =  { ( n506 ) , ( n595 ) }  ;
assign n597 =  { ( n489 ) , ( n596 ) }  ;
assign n598 =  { ( n472 ) , ( n597 ) }  ;
assign n599 =  { ( n455 ) , ( n598 ) }  ;
assign n600 =  ( n438 ) ? ( n599 ) : ( stencil_stream_buff_0 ) ;
assign n601 =  ( n37 ) ? ( stencil_stream_buff_0 ) : ( stencil_stream_buff_0 ) ;
assign n602 =  ( n32 ) ? ( stencil_stream_buff_0 ) : ( n601 ) ;
assign n603 =  ( n25 ) ? ( n600 ) : ( n602 ) ;
assign n604 =  ( n18 ) ? ( stencil_stream_buff_0 ) : ( n603 ) ;
assign n605 =  ( n9 ) ? ( stencil_stream_buff_0 ) : ( n604 ) ;
assign n606 =  ( n4 ) ? ( stencil_stream_buff_0 ) : ( n605 ) ;
assign n607 =  ( n37 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_1 ) ;
assign n608 =  ( n32 ) ? ( stencil_stream_buff_1 ) : ( n607 ) ;
assign n609 =  ( n25 ) ? ( stencil_stream_buff_0 ) : ( n608 ) ;
assign n610 =  ( n18 ) ? ( stencil_stream_buff_1 ) : ( n609 ) ;
assign n611 =  ( n9 ) ? ( stencil_stream_buff_1 ) : ( n610 ) ;
assign n612 =  ( n4 ) ? ( stencil_stream_buff_1 ) : ( n611 ) ;
assign n613 =  ( n162 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n614 =  ( n23 ) ? ( stencil_stream_empty ) : ( 1'd0 ) ;
assign n615 =  ( n37 ) ? ( stencil_stream_empty ) : ( stencil_stream_empty ) ;
assign n616 =  ( n32 ) ? ( stencil_stream_empty ) : ( n615 ) ;
assign n617 =  ( n25 ) ? ( n614 ) : ( n616 ) ;
assign n618 =  ( n18 ) ? ( n613 ) : ( n617 ) ;
assign n619 =  ( n9 ) ? ( stencil_stream_empty ) : ( n618 ) ;
assign n620 =  ( n4 ) ? ( stencil_stream_empty ) : ( n619 ) ;
assign n621 =  ( n14 ) ? ( 1'd0 ) : ( 1'd0 ) ;
assign n622 =  ( stencil_stream_empty ) == ( 1'd1 )  ;
assign n623 =  ( n622 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n624 =  ( n23 ) ? ( stencil_stream_full ) : ( n623 ) ;
assign n625 =  ( n37 ) ? ( stencil_stream_full ) : ( stencil_stream_full ) ;
assign n626 =  ( n32 ) ? ( stencil_stream_full ) : ( n625 ) ;
assign n627 =  ( n25 ) ? ( n624 ) : ( n626 ) ;
assign n628 =  ( n18 ) ? ( n621 ) : ( n627 ) ;
assign n629 =  ( n9 ) ? ( stencil_stream_full ) : ( n628 ) ;
assign n630 =  ( n4 ) ? ( stencil_stream_full ) : ( n629 ) ;
assign n631 = ~ ( n4 ) ;
assign n632 = ~ ( n9 ) ;
assign n633 =  ( n631 ) & ( n632 )  ;
assign n634 = ~ ( n18 ) ;
assign n635 =  ( n633 ) & ( n634 )  ;
assign n636 = ~ ( n25 ) ;
assign n637 =  ( n635 ) & ( n636 )  ;
assign n638 = ~ ( n32 ) ;
assign n639 =  ( n637 ) & ( n638 )  ;
assign n640 = ~ ( n37 ) ;
assign n641 =  ( n639 ) & ( n640 )  ;
assign n642 =  ( n639 ) & ( n37 )  ;
assign n643 =  ( n637 ) & ( n32 )  ;
assign n644 = ~ ( n328 ) ;
assign n645 =  ( n643 ) & ( n644 )  ;
assign n646 =  ( n643 ) & ( n328 )  ;
assign n647 =  ( n635 ) & ( n25 )  ;
assign n648 =  ( n633 ) & ( n18 )  ;
assign n649 =  ( n631 ) & ( n9 )  ;
assign LB2D_proc_0_addr0 = n646 ? (LB2D_proc_x) : (0);
assign LB2D_proc_0_data0 = n646 ? (n327) : (LB2D_proc_0[0]);
assign n650 = ~ ( n330 ) ;
assign n651 =  ( n643 ) & ( n650 )  ;
assign n652 =  ( n643 ) & ( n330 )  ;
assign LB2D_proc_1_addr0 = n652 ? (LB2D_proc_x) : (0);
assign LB2D_proc_1_data0 = n652 ? (n327) : (LB2D_proc_1[0]);
assign n653 = ~ ( n332 ) ;
assign n654 =  ( n643 ) & ( n653 )  ;
assign n655 =  ( n643 ) & ( n332 )  ;
assign LB2D_proc_2_addr0 = n655 ? (LB2D_proc_x) : (0);
assign LB2D_proc_2_data0 = n655 ? (n327) : (LB2D_proc_2[0]);
assign n656 = ~ ( n334 ) ;
assign n657 =  ( n643 ) & ( n656 )  ;
assign n658 =  ( n643 ) & ( n334 )  ;
assign LB2D_proc_3_addr0 = n658 ? (LB2D_proc_x) : (0);
assign LB2D_proc_3_data0 = n658 ? (n327) : (LB2D_proc_3[0]);
assign n659 = ~ ( n336 ) ;
assign n660 =  ( n643 ) & ( n659 )  ;
assign n661 =  ( n643 ) & ( n336 )  ;
assign LB2D_proc_4_addr0 = n661 ? (LB2D_proc_x) : (0);
assign LB2D_proc_4_data0 = n661 ? (n327) : (LB2D_proc_4[0]);
assign n662 = ~ ( n338 ) ;
assign n663 =  ( n643 ) & ( n662 )  ;
assign n664 =  ( n643 ) & ( n338 )  ;
assign LB2D_proc_5_addr0 = n664 ? (LB2D_proc_x) : (0);
assign LB2D_proc_5_data0 = n664 ? (n327) : (LB2D_proc_5[0]);
assign n665 = ~ ( n340 ) ;
assign n666 =  ( n643 ) & ( n665 )  ;
assign n667 =  ( n643 ) & ( n340 )  ;
assign LB2D_proc_6_addr0 = n667 ? (LB2D_proc_x) : (0);
assign LB2D_proc_6_data0 = n667 ? (n327) : (LB2D_proc_6[0]);
assign n668 =  ( LB2D_proc_w ) == ( 64'd7 )  ;
assign n669 = ~ ( n668 ) ;
assign n670 =  ( n643 ) & ( n669 )  ;
assign n671 =  ( n643 ) & ( n668 )  ;
assign LB2D_proc_7_addr0 = n671 ? (LB2D_proc_x) : (0);
assign LB2D_proc_7_data0 = n671 ? (n327) : (LB2D_proc_7[0]);
function [7:0] gb_fun ;
input [647:0] arg0;
    begin
//TODO: Add the specific function HERE.    end
endfunction

always @(posedge clk) begin
   if(rst) begin
       LB1D_buff <= LB1D_buff;
       LB1D_in <= LB1D_in;
       LB1D_it_1 <= LB1D_it_1;
       LB1D_p_cnt <= LB1D_p_cnt;
       LB2D_proc_w <= LB2D_proc_w;
       LB2D_proc_x <= LB2D_proc_x;
       LB2D_proc_y <= LB2D_proc_y;
       LB2D_shift_0 <= LB2D_shift_0;
       LB2D_shift_1 <= LB2D_shift_1;
       LB2D_shift_2 <= LB2D_shift_2;
       LB2D_shift_3 <= LB2D_shift_3;
       LB2D_shift_4 <= LB2D_shift_4;
       LB2D_shift_5 <= LB2D_shift_5;
       LB2D_shift_6 <= LB2D_shift_6;
       LB2D_shift_7 <= LB2D_shift_7;
       LB2D_shift_x <= LB2D_shift_x;
       LB2D_shift_y <= LB2D_shift_y;
       arg_0_TDATA <= arg_0_TDATA;
       arg_0_TVALID <= arg_0_TVALID;
       arg_1_TREADY <= arg_1_TREADY;
       gb_exit_it_1 <= gb_exit_it_1;
       gb_exit_it_2 <= gb_exit_it_2;
       gb_exit_it_3 <= gb_exit_it_3;
       gb_exit_it_4 <= gb_exit_it_4;
       gb_exit_it_5 <= gb_exit_it_5;
       gb_exit_it_6 <= gb_exit_it_6;
       gb_exit_it_7 <= gb_exit_it_7;
       gb_exit_it_8 <= gb_exit_it_8;
       gb_p_cnt <= gb_p_cnt;
       gb_pp_it_1 <= gb_pp_it_1;
       gb_pp_it_2 <= gb_pp_it_2;
       gb_pp_it_3 <= gb_pp_it_3;
       gb_pp_it_4 <= gb_pp_it_4;
       gb_pp_it_5 <= gb_pp_it_5;
       gb_pp_it_6 <= gb_pp_it_6;
       gb_pp_it_7 <= gb_pp_it_7;
       gb_pp_it_8 <= gb_pp_it_8;
       gb_pp_it_9 <= gb_pp_it_9;
       in_stream_buff_0 <= in_stream_buff_0;
       in_stream_buff_1 <= in_stream_buff_1;
       in_stream_empty <= in_stream_empty;
       in_stream_full <= in_stream_full;
       slice_stream_buff_0 <= slice_stream_buff_0;
       slice_stream_buff_1 <= slice_stream_buff_1;
       slice_stream_empty <= slice_stream_empty;
       slice_stream_full <= slice_stream_full;
       stencil_stream_buff_0 <= stencil_stream_buff_0;
       stencil_stream_buff_1 <= stencil_stream_buff_1;
       stencil_stream_empty <= stencil_stream_empty;
       stencil_stream_full <= stencil_stream_full;
   end
   else if(step) begin
       LB1D_buff <= n43;
       LB1D_in <= n49;
       LB1D_it_1 <= n52;
       LB1D_p_cnt <= n63;
       LB2D_proc_w <= n74;
       LB2D_proc_x <= n85;
       LB2D_proc_y <= n93;
       LB2D_shift_0 <= n101;
       LB2D_shift_1 <= n107;
       LB2D_shift_2 <= n113;
       LB2D_shift_3 <= n119;
       LB2D_shift_4 <= n125;
       LB2D_shift_5 <= n131;
       LB2D_shift_6 <= n137;
       LB2D_shift_7 <= n143;
       LB2D_shift_x <= n150;
       LB2D_shift_y <= n161;
       arg_0_TDATA <= n170;
       arg_0_TVALID <= n178;
       arg_1_TREADY <= n185;
       gb_exit_it_1 <= n194;
       gb_exit_it_2 <= n200;
       gb_exit_it_3 <= n206;
       gb_exit_it_4 <= n212;
       gb_exit_it_5 <= n218;
       gb_exit_it_6 <= n224;
       gb_exit_it_7 <= n230;
       gb_exit_it_8 <= n236;
       gb_p_cnt <= n244;
       gb_pp_it_1 <= n250;
       gb_pp_it_2 <= n256;
       gb_pp_it_3 <= n262;
       gb_pp_it_4 <= n268;
       gb_pp_it_5 <= n274;
       gb_pp_it_6 <= n280;
       gb_pp_it_7 <= n286;
       gb_pp_it_8 <= n292;
       gb_pp_it_9 <= n298;
       in_stream_buff_0 <= n304;
       in_stream_buff_1 <= n310;
       in_stream_empty <= n318;
       in_stream_full <= n326;
       slice_stream_buff_0 <= n413;
       slice_stream_buff_1 <= n420;
       slice_stream_empty <= n428;
       slice_stream_full <= n437;
       stencil_stream_buff_0 <= n606;
       stencil_stream_buff_1 <= n612;
       stencil_stream_empty <= n620;
       stencil_stream_full <= n630;
       LB2D_proc_0 [ LB2D_proc_0_addr0 ] <= LB2D_proc_0_data0;
       LB2D_proc_1 [ LB2D_proc_1_addr0 ] <= LB2D_proc_1_data0;
       LB2D_proc_2 [ LB2D_proc_2_addr0 ] <= LB2D_proc_2_data0;
       LB2D_proc_3 [ LB2D_proc_3_addr0 ] <= LB2D_proc_3_data0;
       LB2D_proc_4 [ LB2D_proc_4_addr0 ] <= LB2D_proc_4_data0;
       LB2D_proc_5 [ LB2D_proc_5_addr0 ] <= LB2D_proc_5_data0;
       LB2D_proc_6 [ LB2D_proc_6_addr0 ] <= LB2D_proc_6_data0;
       LB2D_proc_7 [ LB2D_proc_7_addr0 ] <= LB2D_proc_7_data0;
   end
end
endmodule
