module GB(
arg_0_TREADY,
arg_1_TDATA,
arg_1_TVALID,
RAM_w,
RAM_x,
RAM_y,
arg_0_TDATA,
arg_0_TVALID,
arg_1_TREADY,
proc_in,
stencil_0,
stencil_1,
stencil_2,
stencil_3,
stencil_4,
stencil_5,
stencil_6,
stencil_7,
stencil_8,
clk,rst,
step
);
input            arg_0_TREADY;
input      [7:0] arg_1_TDATA;
input            arg_1_TVALID;
input clk;
input rst;
input step;
output      [2:0] RAM_w;
output      [8:0] RAM_x;
output      [9:0] RAM_y;
output      [7:0] arg_0_TDATA;
output            arg_0_TVALID;
output            arg_1_TREADY;
output    [647:0] proc_in;
output     [71:0] stencil_0;
output     [71:0] stencil_1;
output     [71:0] stencil_2;
output     [71:0] stencil_3;
output     [71:0] stencil_4;
output     [71:0] stencil_5;
output     [71:0] stencil_6;
output     [71:0] stencil_7;
output     [71:0] stencil_8;
reg      [2:0] RAM_w;
reg      [8:0] RAM_x;
reg      [9:0] RAM_y;
reg      [7:0] arg_0_TDATA;
reg            arg_0_TVALID;
reg            arg_1_TREADY;
reg    [647:0] proc_in;
reg     [71:0] stencil_0;
reg     [71:0] stencil_1;
reg     [71:0] stencil_2;
reg     [71:0] stencil_3;
reg     [71:0] stencil_4;
reg     [71:0] stencil_5;
reg     [71:0] stencil_6;
reg     [71:0] stencil_7;
reg     [71:0] stencil_8;
wire            arg_0_TREADY;
wire      [7:0] arg_1_TDATA;
wire            arg_1_TVALID;
wire            n0;
wire            n1;
wire            n2;
wire            n3;
wire      [2:0] n4;
wire      [2:0] n5;
wire      [2:0] n6;
wire      [2:0] n7;
wire      [2:0] n8;
wire      [8:0] n9;
wire      [8:0] n10;
wire      [8:0] n11;
wire      [8:0] n12;
wire            n13;
wire      [9:0] n14;
wire      [9:0] n15;
wire      [9:0] n16;
wire      [9:0] n17;
wire      [9:0] n18;
wire            n19;
wire      [7:0] n20;
wire      [7:0] n21;
wire      [7:0] n22;
wire      [7:0] n23;
wire      [7:0] n24;
wire      [7:0] n25;
wire      [7:0] n26;
wire      [7:0] n27;
wire      [7:0] n28;
wire     [15:0] n29;
wire     [23:0] n30;
wire     [31:0] n31;
wire     [39:0] n32;
wire     [47:0] n33;
wire     [55:0] n34;
wire     [63:0] n35;
wire     [71:0] n36;
wire      [7:0] n37;
wire      [7:0] n38;
wire      [7:0] n39;
wire      [7:0] n40;
wire      [7:0] n41;
wire      [7:0] n42;
wire      [7:0] n43;
wire      [7:0] n44;
wire      [7:0] n45;
wire     [15:0] n46;
wire     [23:0] n47;
wire     [31:0] n48;
wire     [39:0] n49;
wire     [47:0] n50;
wire     [55:0] n51;
wire     [63:0] n52;
wire     [71:0] n53;
wire      [7:0] n54;
wire      [7:0] n55;
wire      [7:0] n56;
wire      [7:0] n57;
wire      [7:0] n58;
wire      [7:0] n59;
wire      [7:0] n60;
wire      [7:0] n61;
wire      [7:0] n62;
wire     [15:0] n63;
wire     [23:0] n64;
wire     [31:0] n65;
wire     [39:0] n66;
wire     [47:0] n67;
wire     [55:0] n68;
wire     [63:0] n69;
wire     [71:0] n70;
wire      [7:0] n71;
wire      [7:0] n72;
wire      [7:0] n73;
wire      [7:0] n74;
wire      [7:0] n75;
wire      [7:0] n76;
wire      [7:0] n77;
wire      [7:0] n78;
wire      [7:0] n79;
wire     [15:0] n80;
wire     [23:0] n81;
wire     [31:0] n82;
wire     [39:0] n83;
wire     [47:0] n84;
wire     [55:0] n85;
wire     [63:0] n86;
wire     [71:0] n87;
wire      [7:0] n88;
wire      [7:0] n89;
wire      [7:0] n90;
wire      [7:0] n91;
wire      [7:0] n92;
wire      [7:0] n93;
wire      [7:0] n94;
wire      [7:0] n95;
wire      [7:0] n96;
wire     [15:0] n97;
wire     [23:0] n98;
wire     [31:0] n99;
wire     [39:0] n100;
wire     [47:0] n101;
wire     [55:0] n102;
wire     [63:0] n103;
wire     [71:0] n104;
wire      [7:0] n105;
wire      [7:0] n106;
wire      [7:0] n107;
wire      [7:0] n108;
wire      [7:0] n109;
wire      [7:0] n110;
wire      [7:0] n111;
wire      [7:0] n112;
wire      [7:0] n113;
wire     [15:0] n114;
wire     [23:0] n115;
wire     [31:0] n116;
wire     [39:0] n117;
wire     [47:0] n118;
wire     [55:0] n119;
wire     [63:0] n120;
wire     [71:0] n121;
wire      [7:0] n122;
wire      [7:0] n123;
wire      [7:0] n124;
wire      [7:0] n125;
wire      [7:0] n126;
wire      [7:0] n127;
wire      [7:0] n128;
wire      [7:0] n129;
wire      [7:0] n130;
wire     [15:0] n131;
wire     [23:0] n132;
wire     [31:0] n133;
wire     [39:0] n134;
wire     [47:0] n135;
wire     [55:0] n136;
wire     [63:0] n137;
wire     [71:0] n138;
wire      [7:0] n139;
wire      [7:0] n140;
wire      [7:0] n141;
wire      [7:0] n142;
wire      [7:0] n143;
wire      [7:0] n144;
wire      [7:0] n145;
wire      [7:0] n146;
wire      [7:0] n147;
wire     [15:0] n148;
wire     [23:0] n149;
wire     [31:0] n150;
wire     [39:0] n151;
wire     [47:0] n152;
wire     [55:0] n153;
wire     [63:0] n154;
wire     [71:0] n155;
wire      [7:0] n156;
wire      [7:0] n157;
wire      [7:0] n158;
wire      [7:0] n159;
wire      [7:0] n160;
wire      [7:0] n161;
wire      [7:0] n162;
wire      [7:0] n163;
wire      [7:0] n164;
wire     [15:0] n165;
wire     [23:0] n166;
wire     [31:0] n167;
wire     [39:0] n168;
wire     [47:0] n169;
wire     [55:0] n170;
wire     [63:0] n171;
wire     [71:0] n172;
wire    [143:0] n173;
wire    [215:0] n174;
wire    [287:0] n175;
wire    [359:0] n176;
wire    [431:0] n177;
wire    [503:0] n178;
wire    [575:0] n179;
wire    [647:0] n180;
wire    [647:0] n181;
wire      [7:0] n182;
wire      [7:0] n183;
wire      [7:0] n184;
wire            n185;
wire            n186;
wire            n187;
wire            n188;
wire            n189;
wire    [647:0] n190;
wire      [8:0] RAM_0_addr0;
wire      [7:0] RAM_0_data0;
wire            n191;
wire            n192;
wire            n193;
wire            n194;
wire            n195;
wire            n196;
wire            n197;
wire      [8:0] n198;
wire      [8:0] RAM_1_addr0;
wire      [7:0] RAM_1_data0;
wire            n199;
wire            n200;
wire            n201;
wire            n202;
wire      [8:0] RAM_2_addr0;
wire      [7:0] RAM_2_data0;
wire            n203;
wire            n204;
wire            n205;
wire            n206;
wire      [8:0] RAM_3_addr0;
wire      [7:0] RAM_3_data0;
wire            n207;
wire            n208;
wire            n209;
wire            n210;
wire      [8:0] RAM_4_addr0;
wire      [7:0] RAM_4_data0;
wire            n211;
wire            n212;
wire            n213;
wire            n214;
wire      [8:0] RAM_5_addr0;
wire      [7:0] RAM_5_data0;
wire            n215;
wire            n216;
wire            n217;
wire            n218;
wire      [8:0] RAM_6_addr0;
wire      [7:0] RAM_6_data0;
wire            n219;
wire            n220;
wire            n221;
wire            n222;
wire      [8:0] RAM_7_addr0;
wire      [7:0] RAM_7_data0;
wire            n223;
wire            n224;
wire            n225;
reg      [7:0] RAM_0[511:0];
reg      [7:0] RAM_1[511:0];
reg      [7:0] RAM_2[511:0];
reg      [7:0] RAM_3[511:0];
reg      [7:0] RAM_4[511:0];
reg      [7:0] RAM_5[511:0];
reg      [7:0] RAM_6[511:0];
reg      [7:0] RAM_7[511:0];
wire clk;
wire rst;
wire step;
assign n0 =  ( 1'd0 ) & ( arg_0_TREADY )  ;
assign n1 =  ( n0 ) == ( 1'd0 )  ;
assign n2 =  ( RAM_x ) == ( 9'd488 )  ;
assign n3 =  ( RAM_w ) == ( 3'd7 )  ;
assign n4 =  ( RAM_w ) + ( 3'd1 )  ;
assign n5 =  ( n3 ) ? ( 3'd0 ) : ( n4 ) ;
assign n6 =  ( n2 ) ? ( n5 ) : ( RAM_w ) ;
assign n7 =  ( n1 ) ? ( n6 ) : ( RAM_w ) ;
assign n8 =  ( n1 ) ? ( RAM_w ) : ( n7 ) ;
assign n9 =  ( RAM_x ) + ( 9'd1 )  ;
assign n10 =  ( n2 ) ? ( 9'd1 ) : ( n9 ) ;
assign n11 =  ( n1 ) ? ( n10 ) : ( RAM_x ) ;
assign n12 =  ( n1 ) ? ( RAM_x ) : ( n11 ) ;
assign n13 =  ( RAM_y ) == ( 10'd648 )  ;
assign n14 =  ( RAM_y ) + ( 10'd1 )  ;
assign n15 =  ( n13 ) ? ( 10'd0 ) : ( n14 ) ;
assign n16 =  ( n2 ) ? ( n15 ) : ( RAM_y ) ;
assign n17 =  ( n1 ) ? ( n16 ) : ( RAM_y ) ;
assign n18 =  ( n1 ) ? ( RAM_y ) : ( n17 ) ;
assign n19 =  ( RAM_x ) > ( 9'd9 )  ;
assign n20 = stencil_8[71:64] ;
assign n21 = stencil_7[71:64] ;
assign n22 = stencil_6[71:64] ;
assign n23 = stencil_5[71:64] ;
assign n24 = stencil_4[71:64] ;
assign n25 = stencil_3[71:64] ;
assign n26 = stencil_2[71:64] ;
assign n27 = stencil_1[71:64] ;
assign n28 = stencil_0[71:64] ;
assign n29 =  { ( n27 ) , ( n28 ) }  ;
assign n30 =  { ( n26 ) , ( n29 ) }  ;
assign n31 =  { ( n25 ) , ( n30 ) }  ;
assign n32 =  { ( n24 ) , ( n31 ) }  ;
assign n33 =  { ( n23 ) , ( n32 ) }  ;
assign n34 =  { ( n22 ) , ( n33 ) }  ;
assign n35 =  { ( n21 ) , ( n34 ) }  ;
assign n36 =  { ( n20 ) , ( n35 ) }  ;
assign n37 = stencil_8[63:56] ;
assign n38 = stencil_7[63:56] ;
assign n39 = stencil_6[63:56] ;
assign n40 = stencil_5[63:56] ;
assign n41 = stencil_4[63:56] ;
assign n42 = stencil_3[63:56] ;
assign n43 = stencil_2[63:56] ;
assign n44 = stencil_1[63:56] ;
assign n45 = stencil_0[63:56] ;
assign n46 =  { ( n44 ) , ( n45 ) }  ;
assign n47 =  { ( n43 ) , ( n46 ) }  ;
assign n48 =  { ( n42 ) , ( n47 ) }  ;
assign n49 =  { ( n41 ) , ( n48 ) }  ;
assign n50 =  { ( n40 ) , ( n49 ) }  ;
assign n51 =  { ( n39 ) , ( n50 ) }  ;
assign n52 =  { ( n38 ) , ( n51 ) }  ;
assign n53 =  { ( n37 ) , ( n52 ) }  ;
assign n54 = stencil_8[55:48] ;
assign n55 = stencil_7[55:48] ;
assign n56 = stencil_6[55:48] ;
assign n57 = stencil_5[55:48] ;
assign n58 = stencil_4[55:48] ;
assign n59 = stencil_3[55:48] ;
assign n60 = stencil_2[55:48] ;
assign n61 = stencil_1[55:48] ;
assign n62 = stencil_0[55:48] ;
assign n63 =  { ( n61 ) , ( n62 ) }  ;
assign n64 =  { ( n60 ) , ( n63 ) }  ;
assign n65 =  { ( n59 ) , ( n64 ) }  ;
assign n66 =  { ( n58 ) , ( n65 ) }  ;
assign n67 =  { ( n57 ) , ( n66 ) }  ;
assign n68 =  { ( n56 ) , ( n67 ) }  ;
assign n69 =  { ( n55 ) , ( n68 ) }  ;
assign n70 =  { ( n54 ) , ( n69 ) }  ;
assign n71 = stencil_8[47:40] ;
assign n72 = stencil_7[47:40] ;
assign n73 = stencil_6[47:40] ;
assign n74 = stencil_5[47:40] ;
assign n75 = stencil_4[47:40] ;
assign n76 = stencil_3[47:40] ;
assign n77 = stencil_2[47:40] ;
assign n78 = stencil_1[47:40] ;
assign n79 = stencil_0[47:40] ;
assign n80 =  { ( n78 ) , ( n79 ) }  ;
assign n81 =  { ( n77 ) , ( n80 ) }  ;
assign n82 =  { ( n76 ) , ( n81 ) }  ;
assign n83 =  { ( n75 ) , ( n82 ) }  ;
assign n84 =  { ( n74 ) , ( n83 ) }  ;
assign n85 =  { ( n73 ) , ( n84 ) }  ;
assign n86 =  { ( n72 ) , ( n85 ) }  ;
assign n87 =  { ( n71 ) , ( n86 ) }  ;
assign n88 = stencil_8[39:32] ;
assign n89 = stencil_7[39:32] ;
assign n90 = stencil_6[39:32] ;
assign n91 = stencil_5[39:32] ;
assign n92 = stencil_4[39:32] ;
assign n93 = stencil_3[39:32] ;
assign n94 = stencil_2[39:32] ;
assign n95 = stencil_1[39:32] ;
assign n96 = stencil_0[39:32] ;
assign n97 =  { ( n95 ) , ( n96 ) }  ;
assign n98 =  { ( n94 ) , ( n97 ) }  ;
assign n99 =  { ( n93 ) , ( n98 ) }  ;
assign n100 =  { ( n92 ) , ( n99 ) }  ;
assign n101 =  { ( n91 ) , ( n100 ) }  ;
assign n102 =  { ( n90 ) , ( n101 ) }  ;
assign n103 =  { ( n89 ) , ( n102 ) }  ;
assign n104 =  { ( n88 ) , ( n103 ) }  ;
assign n105 = stencil_8[31:24] ;
assign n106 = stencil_7[31:24] ;
assign n107 = stencil_6[31:24] ;
assign n108 = stencil_5[31:24] ;
assign n109 = stencil_4[31:24] ;
assign n110 = stencil_3[31:24] ;
assign n111 = stencil_2[31:24] ;
assign n112 = stencil_1[31:24] ;
assign n113 = stencil_0[31:24] ;
assign n114 =  { ( n112 ) , ( n113 ) }  ;
assign n115 =  { ( n111 ) , ( n114 ) }  ;
assign n116 =  { ( n110 ) , ( n115 ) }  ;
assign n117 =  { ( n109 ) , ( n116 ) }  ;
assign n118 =  { ( n108 ) , ( n117 ) }  ;
assign n119 =  { ( n107 ) , ( n118 ) }  ;
assign n120 =  { ( n106 ) , ( n119 ) }  ;
assign n121 =  { ( n105 ) , ( n120 ) }  ;
assign n122 = stencil_8[23:16] ;
assign n123 = stencil_7[23:16] ;
assign n124 = stencil_6[23:16] ;
assign n125 = stencil_5[23:16] ;
assign n126 = stencil_4[23:16] ;
assign n127 = stencil_3[23:16] ;
assign n128 = stencil_2[23:16] ;
assign n129 = stencil_1[23:16] ;
assign n130 = stencil_0[23:16] ;
assign n131 =  { ( n129 ) , ( n130 ) }  ;
assign n132 =  { ( n128 ) , ( n131 ) }  ;
assign n133 =  { ( n127 ) , ( n132 ) }  ;
assign n134 =  { ( n126 ) , ( n133 ) }  ;
assign n135 =  { ( n125 ) , ( n134 ) }  ;
assign n136 =  { ( n124 ) , ( n135 ) }  ;
assign n137 =  { ( n123 ) , ( n136 ) }  ;
assign n138 =  { ( n122 ) , ( n137 ) }  ;
assign n139 = stencil_8[15:8] ;
assign n140 = stencil_7[15:8] ;
assign n141 = stencil_6[15:8] ;
assign n142 = stencil_5[15:8] ;
assign n143 = stencil_4[15:8] ;
assign n144 = stencil_3[15:8] ;
assign n145 = stencil_2[15:8] ;
assign n146 = stencil_1[15:8] ;
assign n147 = stencil_0[15:8] ;
assign n148 =  { ( n146 ) , ( n147 ) }  ;
assign n149 =  { ( n145 ) , ( n148 ) }  ;
assign n150 =  { ( n144 ) , ( n149 ) }  ;
assign n151 =  { ( n143 ) , ( n150 ) }  ;
assign n152 =  { ( n142 ) , ( n151 ) }  ;
assign n153 =  { ( n141 ) , ( n152 ) }  ;
assign n154 =  { ( n140 ) , ( n153 ) }  ;
assign n155 =  { ( n139 ) , ( n154 ) }  ;
assign n156 = stencil_8[7:0] ;
assign n157 = stencil_7[7:0] ;
assign n158 = stencil_6[7:0] ;
assign n159 = stencil_5[7:0] ;
assign n160 = stencil_4[7:0] ;
assign n161 = stencil_3[7:0] ;
assign n162 = stencil_2[7:0] ;
assign n163 = stencil_1[7:0] ;
assign n164 = stencil_0[7:0] ;
assign n165 =  { ( n163 ) , ( n164 ) }  ;
assign n166 =  { ( n162 ) , ( n165 ) }  ;
assign n167 =  { ( n161 ) , ( n166 ) }  ;
assign n168 =  { ( n160 ) , ( n167 ) }  ;
assign n169 =  { ( n159 ) , ( n168 ) }  ;
assign n170 =  { ( n158 ) , ( n169 ) }  ;
assign n171 =  { ( n157 ) , ( n170 ) }  ;
assign n172 =  { ( n156 ) , ( n171 ) }  ;
assign n173 =  { ( n155 ) , ( n172 ) }  ;
assign n174 =  { ( n138 ) , ( n173 ) }  ;
assign n175 =  { ( n121 ) , ( n174 ) }  ;
assign n176 =  { ( n104 ) , ( n175 ) }  ;
assign n177 =  { ( n87 ) , ( n176 ) }  ;
assign n178 =  { ( n70 ) , ( n177 ) }  ;
assign n179 =  { ( n53 ) , ( n178 ) }  ;
assign n180 =  { ( n36 ) , ( n179 ) }  ;
assign n181 =  ( n19 ) ? ( n180 ) : ( proc_in ) ;
assign n182 = gb_fun(n181) ;
assign n183 =  ( n1 ) ? ( arg_0_TDATA ) : ( arg_0_TDATA ) ;
assign n184 =  ( n1 ) ? ( n182 ) : ( n183 ) ;
assign n185 =  ( n19 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n186 =  ( n1 ) ? ( 1'd0 ) : ( arg_0_TVALID ) ;
assign n187 =  ( n1 ) ? ( n185 ) : ( n186 ) ;
assign n188 =  ( n1 ) ? ( 1'd0 ) : ( arg_1_TREADY ) ;
assign n189 =  ( n1 ) ? ( 1'd1 ) : ( n188 ) ;
assign n190 =  ( n1 ) ? ( n181 ) : ( proc_in ) ;
assign n191 = ~ ( n1 ) ;
assign n192 =  ( n191 ) & ( n191 )  ;
assign n193 =  ( n191 ) & ( n1 )  ;
assign n194 =  ( RAM_w ) == ( 3'd0 )  ;
assign n195 = ~ ( n194 ) ;
assign n196 =  ( n193 ) & ( n195 )  ;
assign n197 =  ( n193 ) & ( n194 )  ;
assign n198 =  ( RAM_x ) - ( 9'd1 )  ;
assign RAM_0_addr0 = n197 ? (n198) : (0);
assign RAM_0_data0 = n197 ? (arg_1_TDATA) : (RAM_0[0]);
assign n199 =  ( RAM_w ) == ( 3'd1 )  ;
assign n200 = ~ ( n199 ) ;
assign n201 =  ( n193 ) & ( n200 )  ;
assign n202 =  ( n193 ) & ( n199 )  ;
assign RAM_1_addr0 = n202 ? (n198) : (0);
assign RAM_1_data0 = n202 ? (arg_1_TDATA) : (RAM_1[0]);
assign n203 =  ( RAM_w ) == ( 3'd2 )  ;
assign n204 = ~ ( n203 ) ;
assign n205 =  ( n193 ) & ( n204 )  ;
assign n206 =  ( n193 ) & ( n203 )  ;
assign RAM_2_addr0 = n206 ? (n198) : (0);
assign RAM_2_data0 = n206 ? (arg_1_TDATA) : (RAM_2[0]);
assign n207 =  ( RAM_w ) == ( 3'd3 )  ;
assign n208 = ~ ( n207 ) ;
assign n209 =  ( n193 ) & ( n208 )  ;
assign n210 =  ( n193 ) & ( n207 )  ;
assign RAM_3_addr0 = n210 ? (n198) : (0);
assign RAM_3_data0 = n210 ? (arg_1_TDATA) : (RAM_3[0]);
assign n211 =  ( RAM_w ) == ( 3'd4 )  ;
assign n212 = ~ ( n211 ) ;
assign n213 =  ( n193 ) & ( n212 )  ;
assign n214 =  ( n193 ) & ( n211 )  ;
assign RAM_4_addr0 = n214 ? (n198) : (0);
assign RAM_4_data0 = n214 ? (arg_1_TDATA) : (RAM_4[0]);
assign n215 =  ( RAM_w ) == ( 3'd5 )  ;
assign n216 = ~ ( n215 ) ;
assign n217 =  ( n193 ) & ( n216 )  ;
assign n218 =  ( n193 ) & ( n215 )  ;
assign RAM_5_addr0 = n218 ? (n198) : (0);
assign RAM_5_data0 = n218 ? (arg_1_TDATA) : (RAM_5[0]);
assign n219 =  ( RAM_w ) == ( 3'd6 )  ;
assign n220 = ~ ( n219 ) ;
assign n221 =  ( n193 ) & ( n220 )  ;
assign n222 =  ( n193 ) & ( n219 )  ;
assign RAM_6_addr0 = n222 ? (n198) : (0);
assign RAM_6_data0 = n222 ? (arg_1_TDATA) : (RAM_6[0]);
assign n223 = ~ ( n3 ) ;
assign n224 =  ( n193 ) & ( n223 )  ;
assign n225 =  ( n193 ) & ( n3 )  ;
assign RAM_7_addr0 = n225 ? (n198) : (0);
assign RAM_7_data0 = n225 ? (arg_1_TDATA) : (RAM_7[0]);
function [7:0] gb_fun ;
input [647:0] arg0;
    begin
//TODO: Add the specific function HERE.    end
endfunction

always @(posedge clk) begin
   if(rst) begin
       RAM_w <= RAM_w;
       RAM_x <= RAM_x;
       RAM_y <= RAM_y;
       arg_0_TDATA <= arg_0_TDATA;
       arg_0_TVALID <= arg_0_TVALID;
       arg_1_TREADY <= arg_1_TREADY;
       proc_in <= proc_in;
       stencil_0 <= stencil_0;
       stencil_1 <= stencil_1;
       stencil_2 <= stencil_2;
       stencil_3 <= stencil_3;
       stencil_4 <= stencil_4;
       stencil_5 <= stencil_5;
       stencil_6 <= stencil_6;
       stencil_7 <= stencil_7;
       stencil_8 <= stencil_8;
   end
   else if(step) begin
       RAM_w <= n8;
       RAM_x <= n12;
       RAM_y <= n18;
       arg_0_TDATA <= n184;
       arg_0_TVALID <= n187;
       arg_1_TREADY <= n189;
       proc_in <= n190;
       RAM_0 [ RAM_0_addr0 ] <= RAM_0_data0;
       RAM_1 [ RAM_1_addr0 ] <= RAM_1_data0;
       RAM_2 [ RAM_2_addr0 ] <= RAM_2_data0;
       RAM_3 [ RAM_3_addr0 ] <= RAM_3_data0;
       RAM_4 [ RAM_4_addr0 ] <= RAM_4_data0;
       RAM_5 [ RAM_5_addr0 ] <= RAM_5_data0;
       RAM_6 [ RAM_6_addr0 ] <= RAM_6_data0;
       RAM_7 [ RAM_7_addr0 ] <= RAM_7_data0;
   end
end
endmodule
