module GB(
arg_0_TREADY,
arg_1_TDATA,
arg_1_TVALID,
LB1D_buff,
LB1D_it_1,
LB1D_p_cnt,
LB2D_proc_w,
LB2D_proc_x,
LB2D_proc_y,
LB2D_shift_0,
LB2D_shift_1,
LB2D_shift_2,
LB2D_shift_3,
LB2D_shift_4,
LB2D_shift_5,
LB2D_shift_6,
LB2D_shift_7,
LB2D_shift_x,
LB2D_shift_y,
arg_0_TDATA,
arg_0_TVALID,
arg_1_TREADY,
gb_exit_it_1,
gb_exit_it_2,
gb_exit_it_3,
gb_exit_it_4,
gb_exit_it_5,
gb_exit_it_6,
gb_exit_it_7,
gb_exit_it_8,
gb_p_cnt,
gb_pp_it_1,
gb_pp_it_2,
gb_pp_it_3,
gb_pp_it_4,
gb_pp_it_5,
gb_pp_it_6,
gb_pp_it_7,
gb_pp_it_8,
gb_pp_it_9,
in_stream_buff_0,
in_stream_buff_1,
in_stream_empty,
in_stream_full,
slice_stream_buff_0,
slice_stream_buff_1,
slice_stream_empty,
slice_stream_full,
stencil_stream_buff_0,
stencil_stream_buff_1,
stencil_stream_empty,
stencil_stream_full,
clk,rst,
step
);
input            arg_0_TREADY;
input      [7:0] arg_1_TDATA;
input            arg_1_TVALID;
input clk;
input rst;
input step;
output      [7:0] LB1D_buff;
output            LB1D_it_1;
output     [18:0] LB1D_p_cnt;
output     [63:0] LB2D_proc_w;
output      [8:0] LB2D_proc_x;
output      [9:0] LB2D_proc_y;
output     [71:0] LB2D_shift_0;
output     [71:0] LB2D_shift_1;
output     [71:0] LB2D_shift_2;
output     [71:0] LB2D_shift_3;
output     [71:0] LB2D_shift_4;
output     [71:0] LB2D_shift_5;
output     [71:0] LB2D_shift_6;
output     [71:0] LB2D_shift_7;
output      [8:0] LB2D_shift_x;
output      [9:0] LB2D_shift_y;
output      [7:0] arg_0_TDATA;
output            arg_0_TVALID;
output            arg_1_TREADY;
output            gb_exit_it_1;
output            gb_exit_it_2;
output            gb_exit_it_3;
output            gb_exit_it_4;
output            gb_exit_it_5;
output            gb_exit_it_6;
output            gb_exit_it_7;
output            gb_exit_it_8;
output     [18:0] gb_p_cnt;
output            gb_pp_it_1;
output            gb_pp_it_2;
output            gb_pp_it_3;
output            gb_pp_it_4;
output            gb_pp_it_5;
output            gb_pp_it_6;
output            gb_pp_it_7;
output            gb_pp_it_8;
output            gb_pp_it_9;
output      [7:0] in_stream_buff_0;
output      [7:0] in_stream_buff_1;
output            in_stream_empty;
output            in_stream_full;
output     [71:0] slice_stream_buff_0;
output     [71:0] slice_stream_buff_1;
output            slice_stream_empty;
output            slice_stream_full;
output    [647:0] stencil_stream_buff_0;
output    [647:0] stencil_stream_buff_1;
output            stencil_stream_empty;
output            stencil_stream_full;
reg      [7:0] LB1D_buff;
reg            LB1D_it_1;
reg     [18:0] LB1D_p_cnt;
reg     [63:0] LB2D_proc_w;
reg      [8:0] LB2D_proc_x;
reg      [9:0] LB2D_proc_y;
reg     [71:0] LB2D_shift_0;
reg     [71:0] LB2D_shift_1;
reg     [71:0] LB2D_shift_2;
reg     [71:0] LB2D_shift_3;
reg     [71:0] LB2D_shift_4;
reg     [71:0] LB2D_shift_5;
reg     [71:0] LB2D_shift_6;
reg     [71:0] LB2D_shift_7;
reg      [8:0] LB2D_shift_x;
reg      [9:0] LB2D_shift_y;
reg      [7:0] arg_0_TDATA;
reg            arg_0_TVALID;
reg            arg_1_TREADY;
reg            gb_exit_it_1;
reg            gb_exit_it_2;
reg            gb_exit_it_3;
reg            gb_exit_it_4;
reg            gb_exit_it_5;
reg            gb_exit_it_6;
reg            gb_exit_it_7;
reg            gb_exit_it_8;
reg     [18:0] gb_p_cnt;
reg            gb_pp_it_1;
reg            gb_pp_it_2;
reg            gb_pp_it_3;
reg            gb_pp_it_4;
reg            gb_pp_it_5;
reg            gb_pp_it_6;
reg            gb_pp_it_7;
reg            gb_pp_it_8;
reg            gb_pp_it_9;
reg      [7:0] in_stream_buff_0;
reg      [7:0] in_stream_buff_1;
reg            in_stream_empty;
reg            in_stream_full;
reg     [71:0] slice_stream_buff_0;
reg     [71:0] slice_stream_buff_1;
reg            slice_stream_empty;
reg            slice_stream_full;
reg    [647:0] stencil_stream_buff_0;
reg    [647:0] stencil_stream_buff_1;
reg            stencil_stream_empty;
reg            stencil_stream_full;
wire            arg_0_TREADY;
wire      [7:0] arg_1_TDATA;
wire            arg_1_TVALID;
wire            n0;
wire            n1;
wire            n2;
wire            n3;
wire            n4;
wire            n5;
wire            n6;
wire            n7;
wire            n8;
wire            n9;
wire            n10;
wire            n11;
wire            n12;
wire            n13;
wire            n14;
wire            n15;
wire            n16;
wire            n17;
wire            n18;
wire            n19;
wire            n20;
wire            n21;
wire            n22;
wire            n23;
wire            n24;
wire            n25;
wire            n26;
wire            n27;
wire            n28;
wire            n29;
wire            n30;
wire            n31;
wire            n32;
wire            n33;
wire            n34;
wire            n35;
wire            n36;
wire            n37;
wire      [7:0] n38;
wire      [7:0] n39;
wire      [7:0] n40;
wire      [7:0] n41;
wire      [7:0] n42;
wire      [7:0] n43;
wire            n44;
wire            n45;
wire            n46;
wire     [18:0] n47;
wire     [18:0] n48;
wire     [18:0] n49;
wire     [18:0] n50;
wire     [18:0] n51;
wire     [18:0] n52;
wire     [18:0] n53;
wire            n54;
wire            n55;
wire     [63:0] n56;
wire     [63:0] n57;
wire     [63:0] n58;
wire     [63:0] n59;
wire     [63:0] n60;
wire     [63:0] n61;
wire     [63:0] n62;
wire     [63:0] n63;
wire     [63:0] n64;
wire            n65;
wire            n66;
wire            n67;
wire      [8:0] n68;
wire      [8:0] n69;
wire      [8:0] n70;
wire      [8:0] n71;
wire      [8:0] n72;
wire      [8:0] n73;
wire      [8:0] n74;
wire      [8:0] n75;
wire            n76;
wire      [9:0] n77;
wire      [9:0] n78;
wire      [9:0] n79;
wire      [9:0] n80;
wire      [9:0] n81;
wire      [9:0] n82;
wire      [9:0] n83;
wire            n84;
wire     [71:0] n85;
wire     [71:0] n86;
wire     [71:0] n87;
wire     [71:0] n88;
wire     [71:0] n89;
wire     [71:0] n90;
wire     [71:0] n91;
wire     [71:0] n92;
wire     [71:0] n93;
wire     [71:0] n94;
wire     [71:0] n95;
wire     [71:0] n96;
wire     [71:0] n97;
wire     [71:0] n98;
wire     [71:0] n99;
wire     [71:0] n100;
wire     [71:0] n101;
wire     [71:0] n102;
wire     [71:0] n103;
wire     [71:0] n104;
wire     [71:0] n105;
wire     [71:0] n106;
wire     [71:0] n107;
wire     [71:0] n108;
wire     [71:0] n109;
wire     [71:0] n110;
wire     [71:0] n111;
wire     [71:0] n112;
wire     [71:0] n113;
wire     [71:0] n114;
wire     [71:0] n115;
wire     [71:0] n116;
wire     [71:0] n117;
wire     [71:0] n118;
wire     [71:0] n119;
wire     [71:0] n120;
wire     [71:0] n121;
wire     [71:0] n122;
wire     [71:0] n123;
wire     [71:0] n124;
wire     [71:0] n125;
wire     [71:0] n126;
wire     [71:0] n127;
wire     [71:0] n128;
wire     [71:0] n129;
wire     [71:0] n130;
wire     [71:0] n131;
wire     [71:0] n132;
wire     [71:0] n133;
wire            n134;
wire      [8:0] n135;
wire      [8:0] n136;
wire      [8:0] n137;
wire      [8:0] n138;
wire      [8:0] n139;
wire      [8:0] n140;
wire      [8:0] n141;
wire      [8:0] n142;
wire            n143;
wire      [9:0] n144;
wire      [9:0] n145;
wire      [9:0] n146;
wire      [9:0] n147;
wire      [9:0] n148;
wire      [9:0] n149;
wire      [9:0] n150;
wire      [9:0] n151;
wire      [9:0] n152;
wire            n153;
wire    [647:0] n154;
wire      [7:0] n155;
wire      [7:0] n156;
wire      [7:0] n157;
wire      [7:0] n158;
wire      [7:0] n159;
wire      [7:0] n160;
wire      [7:0] n161;
wire            n162;
wire            n163;
wire            n164;
wire            n165;
wire            n166;
wire            n167;
wire            n168;
wire            n169;
wire            n170;
wire            n171;
wire            n172;
wire            n173;
wire            n174;
wire            n175;
wire     [18:0] n176;
wire            n177;
wire            n178;
wire            n179;
wire            n180;
wire            n181;
wire            n182;
wire            n183;
wire            n184;
wire            n185;
wire            n186;
wire            n187;
wire            n188;
wire            n189;
wire            n190;
wire            n191;
wire            n192;
wire            n193;
wire            n194;
wire            n195;
wire            n196;
wire            n197;
wire            n198;
wire            n199;
wire            n200;
wire            n201;
wire            n202;
wire            n203;
wire            n204;
wire            n205;
wire            n206;
wire            n207;
wire            n208;
wire            n209;
wire            n210;
wire            n211;
wire            n212;
wire            n213;
wire            n214;
wire            n215;
wire            n216;
wire            n217;
wire            n218;
wire            n219;
wire            n220;
wire            n221;
wire            n222;
wire            n223;
wire            n224;
wire            n225;
wire            n226;
wire            n227;
wire     [18:0] n228;
wire     [18:0] n229;
wire     [18:0] n230;
wire     [18:0] n231;
wire     [18:0] n232;
wire     [18:0] n233;
wire     [18:0] n234;
wire            n235;
wire            n236;
wire            n237;
wire            n238;
wire            n239;
wire            n240;
wire            n241;
wire            n242;
wire            n243;
wire            n244;
wire            n245;
wire            n246;
wire            n247;
wire            n248;
wire            n249;
wire            n250;
wire            n251;
wire            n252;
wire            n253;
wire            n254;
wire            n255;
wire            n256;
wire            n257;
wire            n258;
wire            n259;
wire            n260;
wire            n261;
wire            n262;
wire            n263;
wire            n264;
wire            n265;
wire            n266;
wire            n267;
wire            n268;
wire            n269;
wire            n270;
wire            n271;
wire            n272;
wire            n273;
wire            n274;
wire            n275;
wire            n276;
wire            n277;
wire            n278;
wire            n279;
wire            n280;
wire            n281;
wire            n282;
wire            n283;
wire            n284;
wire            n285;
wire            n286;
wire            n287;
wire            n288;
wire      [7:0] n289;
wire      [7:0] n290;
wire      [7:0] n291;
wire      [7:0] n292;
wire      [7:0] n293;
wire      [7:0] n294;
wire      [7:0] n295;
wire      [7:0] n296;
wire      [7:0] n297;
wire      [7:0] n298;
wire      [7:0] n299;
wire      [7:0] n300;
wire            n301;
wire            n302;
wire            n303;
wire            n304;
wire            n305;
wire            n306;
wire            n307;
wire            n308;
wire            n309;
wire            n310;
wire            n311;
wire            n312;
wire            n313;
wire            n314;
wire            n315;
wire            n316;
wire      [7:0] n317;
wire            n318;
wire      [7:0] n319;
wire            n320;
wire      [7:0] n321;
wire            n322;
wire      [7:0] n323;
wire            n324;
wire      [7:0] n325;
wire            n326;
wire      [7:0] n327;
wire            n328;
wire      [7:0] n329;
wire            n330;
wire      [7:0] n331;
wire      [7:0] n332;
wire      [7:0] n333;
wire      [7:0] n334;
wire      [7:0] n335;
wire      [7:0] n336;
wire      [7:0] n337;
wire      [7:0] n338;
wire      [7:0] n339;
wire      [7:0] n340;
wire      [7:0] n341;
wire      [7:0] n342;
wire      [7:0] n343;
wire      [7:0] n344;
wire      [7:0] n345;
wire      [7:0] n346;
wire      [7:0] n347;
wire      [7:0] n348;
wire      [7:0] n349;
wire      [7:0] n350;
wire      [7:0] n351;
wire      [7:0] n352;
wire      [7:0] n353;
wire      [7:0] n354;
wire      [7:0] n355;
wire      [7:0] n356;
wire      [7:0] n357;
wire      [7:0] n358;
wire      [7:0] n359;
wire      [7:0] n360;
wire      [7:0] n361;
wire      [7:0] n362;
wire      [7:0] n363;
wire      [7:0] n364;
wire      [7:0] n365;
wire      [7:0] n366;
wire      [7:0] n367;
wire      [7:0] n368;
wire      [7:0] n369;
wire      [7:0] n370;
wire      [7:0] n371;
wire      [7:0] n372;
wire      [7:0] n373;
wire      [7:0] n374;
wire      [7:0] n375;
wire      [7:0] n376;
wire      [7:0] n377;
wire      [7:0] n378;
wire      [7:0] n379;
wire      [7:0] n380;
wire      [7:0] n381;
wire      [7:0] n382;
wire      [7:0] n383;
wire      [7:0] n384;
wire      [7:0] n385;
wire      [7:0] n386;
wire      [7:0] n387;
wire      [7:0] n388;
wire     [15:0] n389;
wire     [23:0] n390;
wire     [31:0] n391;
wire     [39:0] n392;
wire     [47:0] n393;
wire     [55:0] n394;
wire     [63:0] n395;
wire     [71:0] n396;
wire     [71:0] n397;
wire     [71:0] n398;
wire     [71:0] n399;
wire     [71:0] n400;
wire     [71:0] n401;
wire     [71:0] n402;
wire     [71:0] n403;
wire     [71:0] n404;
wire     [71:0] n405;
wire     [71:0] n406;
wire     [71:0] n407;
wire     [71:0] n408;
wire     [71:0] n409;
wire     [71:0] n410;
wire            n411;
wire            n412;
wire            n413;
wire            n414;
wire            n415;
wire            n416;
wire            n417;
wire            n418;
wire            n419;
wire            n420;
wire            n421;
wire            n422;
wire            n423;
wire            n424;
wire            n425;
wire            n426;
wire            n427;
wire            n428;
wire      [7:0] n429;
wire      [7:0] n430;
wire      [7:0] n431;
wire      [7:0] n432;
wire      [7:0] n433;
wire      [7:0] n434;
wire      [7:0] n435;
wire      [7:0] n436;
wire      [7:0] n437;
wire     [15:0] n438;
wire     [23:0] n439;
wire     [31:0] n440;
wire     [39:0] n441;
wire     [47:0] n442;
wire     [55:0] n443;
wire     [63:0] n444;
wire     [71:0] n445;
wire      [7:0] n446;
wire      [7:0] n447;
wire      [7:0] n448;
wire      [7:0] n449;
wire      [7:0] n450;
wire      [7:0] n451;
wire      [7:0] n452;
wire      [7:0] n453;
wire      [7:0] n454;
wire     [15:0] n455;
wire     [23:0] n456;
wire     [31:0] n457;
wire     [39:0] n458;
wire     [47:0] n459;
wire     [55:0] n460;
wire     [63:0] n461;
wire     [71:0] n462;
wire      [7:0] n463;
wire      [7:0] n464;
wire      [7:0] n465;
wire      [7:0] n466;
wire      [7:0] n467;
wire      [7:0] n468;
wire      [7:0] n469;
wire      [7:0] n470;
wire      [7:0] n471;
wire     [15:0] n472;
wire     [23:0] n473;
wire     [31:0] n474;
wire     [39:0] n475;
wire     [47:0] n476;
wire     [55:0] n477;
wire     [63:0] n478;
wire     [71:0] n479;
wire      [7:0] n480;
wire      [7:0] n481;
wire      [7:0] n482;
wire      [7:0] n483;
wire      [7:0] n484;
wire      [7:0] n485;
wire      [7:0] n486;
wire      [7:0] n487;
wire      [7:0] n488;
wire     [15:0] n489;
wire     [23:0] n490;
wire     [31:0] n491;
wire     [39:0] n492;
wire     [47:0] n493;
wire     [55:0] n494;
wire     [63:0] n495;
wire     [71:0] n496;
wire      [7:0] n497;
wire      [7:0] n498;
wire      [7:0] n499;
wire      [7:0] n500;
wire      [7:0] n501;
wire      [7:0] n502;
wire      [7:0] n503;
wire      [7:0] n504;
wire      [7:0] n505;
wire     [15:0] n506;
wire     [23:0] n507;
wire     [31:0] n508;
wire     [39:0] n509;
wire     [47:0] n510;
wire     [55:0] n511;
wire     [63:0] n512;
wire     [71:0] n513;
wire      [7:0] n514;
wire      [7:0] n515;
wire      [7:0] n516;
wire      [7:0] n517;
wire      [7:0] n518;
wire      [7:0] n519;
wire      [7:0] n520;
wire      [7:0] n521;
wire      [7:0] n522;
wire     [15:0] n523;
wire     [23:0] n524;
wire     [31:0] n525;
wire     [39:0] n526;
wire     [47:0] n527;
wire     [55:0] n528;
wire     [63:0] n529;
wire     [71:0] n530;
wire      [7:0] n531;
wire      [7:0] n532;
wire      [7:0] n533;
wire      [7:0] n534;
wire      [7:0] n535;
wire      [7:0] n536;
wire      [7:0] n537;
wire      [7:0] n538;
wire      [7:0] n539;
wire     [15:0] n540;
wire     [23:0] n541;
wire     [31:0] n542;
wire     [39:0] n543;
wire     [47:0] n544;
wire     [55:0] n545;
wire     [63:0] n546;
wire     [71:0] n547;
wire      [7:0] n548;
wire      [7:0] n549;
wire      [7:0] n550;
wire      [7:0] n551;
wire      [7:0] n552;
wire      [7:0] n553;
wire      [7:0] n554;
wire      [7:0] n555;
wire      [7:0] n556;
wire     [15:0] n557;
wire     [23:0] n558;
wire     [31:0] n559;
wire     [39:0] n560;
wire     [47:0] n561;
wire     [55:0] n562;
wire     [63:0] n563;
wire     [71:0] n564;
wire      [7:0] n565;
wire      [7:0] n566;
wire      [7:0] n567;
wire      [7:0] n568;
wire      [7:0] n569;
wire      [7:0] n570;
wire      [7:0] n571;
wire      [7:0] n572;
wire      [7:0] n573;
wire     [15:0] n574;
wire     [23:0] n575;
wire     [31:0] n576;
wire     [39:0] n577;
wire     [47:0] n578;
wire     [55:0] n579;
wire     [63:0] n580;
wire     [71:0] n581;
wire    [143:0] n582;
wire    [215:0] n583;
wire    [287:0] n584;
wire    [359:0] n585;
wire    [431:0] n586;
wire    [503:0] n587;
wire    [575:0] n588;
wire    [647:0] n589;
wire    [647:0] n590;
wire    [647:0] n591;
wire    [647:0] n592;
wire    [647:0] n593;
wire    [647:0] n594;
wire    [647:0] n595;
wire    [647:0] n596;
wire    [647:0] n597;
wire    [647:0] n598;
wire    [647:0] n599;
wire    [647:0] n600;
wire    [647:0] n601;
wire    [647:0] n602;
wire            n603;
wire            n604;
wire            n605;
wire            n606;
wire            n607;
wire            n608;
wire            n609;
wire            n610;
wire            n611;
wire            n612;
wire            n613;
wire            n614;
wire            n615;
wire            n616;
wire            n617;
wire            n618;
wire            n619;
wire            n620;
wire      [8:0] LB2D_proc_0_addr0;
wire      [7:0] LB2D_proc_0_data0;
wire            n621;
wire            n622;
wire            n623;
wire            n624;
wire            n625;
wire            n626;
wire            n627;
wire            n628;
wire            n629;
wire            n630;
wire            n631;
wire            n632;
wire            n633;
wire            n634;
wire            n635;
wire            n636;
wire            n637;
wire            n638;
wire            n639;
wire      [8:0] LB2D_proc_1_addr0;
wire      [7:0] LB2D_proc_1_data0;
wire            n640;
wire            n641;
wire            n642;
wire      [8:0] LB2D_proc_2_addr0;
wire      [7:0] LB2D_proc_2_data0;
wire            n643;
wire            n644;
wire            n645;
wire      [8:0] LB2D_proc_3_addr0;
wire      [7:0] LB2D_proc_3_data0;
wire            n646;
wire            n647;
wire            n648;
wire      [8:0] LB2D_proc_4_addr0;
wire      [7:0] LB2D_proc_4_data0;
wire            n649;
wire            n650;
wire            n651;
wire      [8:0] LB2D_proc_5_addr0;
wire      [7:0] LB2D_proc_5_data0;
wire            n652;
wire            n653;
wire            n654;
wire      [8:0] LB2D_proc_6_addr0;
wire      [7:0] LB2D_proc_6_data0;
wire            n655;
wire            n656;
wire            n657;
wire      [8:0] LB2D_proc_7_addr0;
wire      [7:0] LB2D_proc_7_data0;
wire            n658;
wire            n659;
wire            n660;
wire            n661;
reg      [7:0] LB2D_proc_0[511:0];
reg      [7:0] LB2D_proc_1[511:0];
reg      [7:0] LB2D_proc_2[511:0];
reg      [7:0] LB2D_proc_3[511:0];
reg      [7:0] LB2D_proc_4[511:0];
reg      [7:0] LB2D_proc_5[511:0];
reg      [7:0] LB2D_proc_6[511:0];
reg      [7:0] LB2D_proc_7[511:0];
wire clk;
wire rst;
wire step;
assign n0 =  ( arg_0_TREADY ) == ( 1'd1 )  ;
assign n1 =  ( arg_0_TVALID ) == ( 1'd1 )  ;
assign n2 =  ( n0 ) & ( n1 )  ;
assign n3 =  ( arg_1_TVALID ) == ( 1'd0 )  ;
assign n4 =  ( n2 ) & ( n3 )  ;
assign n5 =  ( arg_1_TREADY ) == ( 1'd1 )  ;
assign n6 =  ( arg_1_TVALID ) == ( 1'd1 )  ;
assign n7 =  ( n5 ) & ( n6 )  ;
assign n8 =  ( arg_0_TREADY ) == ( 1'd0 )  ;
assign n9 =  ( n7 ) & ( n8 )  ;
assign n10 =  ( arg_0_TVALID ) == ( 1'd0 )  ;
assign n11 =  ( gb_exit_it_1 ) == ( 1'd0 )  ;
assign n12 =  ( stencil_stream_empty ) == ( 1'd0 )  ;
assign n13 =  ( n11 ) & ( n12 )  ;
assign n14 =  ( gb_exit_it_1 ) == ( 1'd1 )  ;
assign n15 =  ( gb_exit_it_8 ) == ( 1'd0 )  ;
assign n16 =  ( n14 ) & ( n15 )  ;
assign n17 =  ( n13 ) | ( n16 )  ;
assign n18 =  ( n10 ) & ( n17 )  ;
assign n19 =  ( slice_stream_empty ) == ( 1'd0 )  ;
assign n20 =  ( stencil_stream_full ) == ( 1'd0 )  ;
assign n21 =  ( LB2D_shift_x ) < ( 9'd8 )  ;
assign n22 =  ( n20 ) | ( n21 )  ;
assign n23 =  ( n19 ) & ( n22 )  ;
assign n24 =  ( in_stream_empty ) == ( 1'd0 )  ;
assign n25 =  ( LB2D_proc_x ) != ( 9'd488 )  ;
assign n26 =  ( n24 ) & ( n25 )  ;
assign n27 =  ( slice_stream_full ) == ( 1'd0 )  ;
assign n28 =  ( LB2D_proc_y ) < ( 10'd8 )  ;
assign n29 =  ( n27 ) | ( n28 )  ;
assign n30 =  ( n26 ) & ( n29 )  ;
assign n31 =  ( arg_1_TREADY ) == ( 1'd0 )  ;
assign n32 =  ( in_stream_full ) == ( 1'd0 )  ;
assign n33 =  ( n31 ) & ( n32 )  ;
assign n34 =  ( LB1D_p_cnt ) != ( 19'd316224 )  ;
assign n35 =  ( n33 ) & ( n34 )  ;
assign n36 =  ( LB1D_it_1 ) == ( 1'd1 )  ;
assign n37 =  ( n35 ) & ( n36 )  ;
assign n38 =  ( n37 ) ? ( LB1D_buff ) : ( LB1D_buff ) ;
assign n39 =  ( n30 ) ? ( LB1D_buff ) : ( n38 ) ;
assign n40 =  ( n23 ) ? ( LB1D_buff ) : ( n39 ) ;
assign n41 =  ( n18 ) ? ( LB1D_buff ) : ( n40 ) ;
assign n42 =  ( n9 ) ? ( arg_1_TDATA ) : ( n41 ) ;
assign n43 =  ( n4 ) ? ( arg_1_TDATA ) : ( n42 ) ;
assign n44 =  ( LB1D_it_1 ) == ( 1'd0 )  ;
assign n45 =  ( n35 ) & ( n44 )  ;
assign n46 =  ( n45 ) ? ( 1'd1 ) : ( LB1D_it_1 ) ;
assign n47 =  ( LB1D_p_cnt ) + ( 19'd1 )  ;
assign n48 =  ( n37 ) ? ( n47 ) : ( LB1D_p_cnt ) ;
assign n49 =  ( n30 ) ? ( LB1D_p_cnt ) : ( n48 ) ;
assign n50 =  ( n23 ) ? ( LB1D_p_cnt ) : ( n49 ) ;
assign n51 =  ( n18 ) ? ( LB1D_p_cnt ) : ( n50 ) ;
assign n52 =  ( n9 ) ? ( LB1D_p_cnt ) : ( n51 ) ;
assign n53 =  ( n4 ) ? ( LB1D_p_cnt ) : ( n52 ) ;
assign n54 =  ( LB2D_proc_w ) < ( 64'd7 )  ;
assign n55 =  ( LB2D_proc_x ) < ( 9'd488 )  ;
assign n56 =  ( LB2D_proc_w ) + ( 64'd1 )  ;
assign n57 =  ( n55 ) ? ( LB2D_proc_w ) : ( n56 ) ;
assign n58 =  ( n54 ) ? ( n57 ) : ( 64'd0 ) ;
assign n59 =  ( n37 ) ? ( LB2D_proc_w ) : ( LB2D_proc_w ) ;
assign n60 =  ( n30 ) ? ( n58 ) : ( n59 ) ;
assign n61 =  ( n23 ) ? ( LB2D_proc_w ) : ( n60 ) ;
assign n62 =  ( n18 ) ? ( LB2D_proc_w ) : ( n61 ) ;
assign n63 =  ( n9 ) ? ( LB2D_proc_w ) : ( n62 ) ;
assign n64 =  ( n4 ) ? ( LB2D_proc_w ) : ( n63 ) ;
assign n65 =  ( LB2D_proc_x ) == ( 9'd488 )  ;
assign n66 =  ( n24 ) & ( n65 )  ;
assign n67 =  ( n66 ) & ( n29 )  ;
assign n68 =  ( LB2D_proc_x ) + ( 9'd1 )  ;
assign n69 =  ( n37 ) ? ( LB2D_proc_x ) : ( LB2D_proc_x ) ;
assign n70 =  ( n30 ) ? ( n68 ) : ( n69 ) ;
assign n71 =  ( n67 ) ? ( 9'd0 ) : ( n70 ) ;
assign n72 =  ( n23 ) ? ( LB2D_proc_x ) : ( n71 ) ;
assign n73 =  ( n18 ) ? ( LB2D_proc_x ) : ( n72 ) ;
assign n74 =  ( n9 ) ? ( LB2D_proc_x ) : ( n73 ) ;
assign n75 =  ( n4 ) ? ( LB2D_proc_x ) : ( n74 ) ;
assign n76 =  ( LB2D_proc_y ) < ( 10'd488 )  ;
assign n77 =  ( n76 ) ? ( LB2D_proc_y ) : ( 10'd488 ) ;
assign n78 =  ( n37 ) ? ( LB2D_proc_y ) : ( LB2D_proc_y ) ;
assign n79 =  ( n30 ) ? ( n77 ) : ( n78 ) ;
assign n80 =  ( n23 ) ? ( LB2D_proc_y ) : ( n79 ) ;
assign n81 =  ( n18 ) ? ( LB2D_proc_y ) : ( n80 ) ;
assign n82 =  ( n9 ) ? ( LB2D_proc_y ) : ( n81 ) ;
assign n83 =  ( n4 ) ? ( LB2D_proc_y ) : ( n82 ) ;
assign n84 =  ( slice_stream_full ) == ( 1'd1 )  ;
assign n85 =  ( n84 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n86 =  ( n37 ) ? ( LB2D_shift_0 ) : ( LB2D_shift_0 ) ;
assign n87 =  ( n30 ) ? ( LB2D_shift_0 ) : ( n86 ) ;
assign n88 =  ( n23 ) ? ( n85 ) : ( n87 ) ;
assign n89 =  ( n18 ) ? ( LB2D_shift_0 ) : ( n88 ) ;
assign n90 =  ( n9 ) ? ( LB2D_shift_0 ) : ( n89 ) ;
assign n91 =  ( n4 ) ? ( LB2D_shift_0 ) : ( n90 ) ;
assign n92 =  ( n37 ) ? ( LB2D_shift_1 ) : ( LB2D_shift_1 ) ;
assign n93 =  ( n30 ) ? ( LB2D_shift_1 ) : ( n92 ) ;
assign n94 =  ( n23 ) ? ( LB2D_shift_0 ) : ( n93 ) ;
assign n95 =  ( n18 ) ? ( LB2D_shift_1 ) : ( n94 ) ;
assign n96 =  ( n9 ) ? ( LB2D_shift_1 ) : ( n95 ) ;
assign n97 =  ( n4 ) ? ( LB2D_shift_1 ) : ( n96 ) ;
assign n98 =  ( n37 ) ? ( LB2D_shift_2 ) : ( LB2D_shift_2 ) ;
assign n99 =  ( n30 ) ? ( LB2D_shift_2 ) : ( n98 ) ;
assign n100 =  ( n23 ) ? ( LB2D_shift_1 ) : ( n99 ) ;
assign n101 =  ( n18 ) ? ( LB2D_shift_2 ) : ( n100 ) ;
assign n102 =  ( n9 ) ? ( LB2D_shift_2 ) : ( n101 ) ;
assign n103 =  ( n4 ) ? ( LB2D_shift_2 ) : ( n102 ) ;
assign n104 =  ( n37 ) ? ( LB2D_shift_3 ) : ( LB2D_shift_3 ) ;
assign n105 =  ( n30 ) ? ( LB2D_shift_3 ) : ( n104 ) ;
assign n106 =  ( n23 ) ? ( LB2D_shift_2 ) : ( n105 ) ;
assign n107 =  ( n18 ) ? ( LB2D_shift_3 ) : ( n106 ) ;
assign n108 =  ( n9 ) ? ( LB2D_shift_3 ) : ( n107 ) ;
assign n109 =  ( n4 ) ? ( LB2D_shift_3 ) : ( n108 ) ;
assign n110 =  ( n37 ) ? ( LB2D_shift_4 ) : ( LB2D_shift_4 ) ;
assign n111 =  ( n30 ) ? ( LB2D_shift_4 ) : ( n110 ) ;
assign n112 =  ( n23 ) ? ( LB2D_shift_3 ) : ( n111 ) ;
assign n113 =  ( n18 ) ? ( LB2D_shift_4 ) : ( n112 ) ;
assign n114 =  ( n9 ) ? ( LB2D_shift_4 ) : ( n113 ) ;
assign n115 =  ( n4 ) ? ( LB2D_shift_4 ) : ( n114 ) ;
assign n116 =  ( n37 ) ? ( LB2D_shift_5 ) : ( LB2D_shift_5 ) ;
assign n117 =  ( n30 ) ? ( LB2D_shift_5 ) : ( n116 ) ;
assign n118 =  ( n23 ) ? ( LB2D_shift_4 ) : ( n117 ) ;
assign n119 =  ( n18 ) ? ( LB2D_shift_5 ) : ( n118 ) ;
assign n120 =  ( n9 ) ? ( LB2D_shift_5 ) : ( n119 ) ;
assign n121 =  ( n4 ) ? ( LB2D_shift_5 ) : ( n120 ) ;
assign n122 =  ( n37 ) ? ( LB2D_shift_6 ) : ( LB2D_shift_6 ) ;
assign n123 =  ( n30 ) ? ( LB2D_shift_6 ) : ( n122 ) ;
assign n124 =  ( n23 ) ? ( LB2D_shift_5 ) : ( n123 ) ;
assign n125 =  ( n18 ) ? ( LB2D_shift_6 ) : ( n124 ) ;
assign n126 =  ( n9 ) ? ( LB2D_shift_6 ) : ( n125 ) ;
assign n127 =  ( n4 ) ? ( LB2D_shift_6 ) : ( n126 ) ;
assign n128 =  ( n37 ) ? ( LB2D_shift_7 ) : ( LB2D_shift_7 ) ;
assign n129 =  ( n30 ) ? ( LB2D_shift_7 ) : ( n128 ) ;
assign n130 =  ( n23 ) ? ( LB2D_shift_6 ) : ( n129 ) ;
assign n131 =  ( n18 ) ? ( LB2D_shift_7 ) : ( n130 ) ;
assign n132 =  ( n9 ) ? ( LB2D_shift_7 ) : ( n131 ) ;
assign n133 =  ( n4 ) ? ( LB2D_shift_7 ) : ( n132 ) ;
assign n134 =  ( LB2D_shift_x ) < ( 9'd487 )  ;
assign n135 =  ( LB2D_shift_x ) + ( 9'd1 )  ;
assign n136 =  ( n134 ) ? ( n135 ) : ( 9'd0 ) ;
assign n137 =  ( n37 ) ? ( LB2D_shift_x ) : ( LB2D_shift_x ) ;
assign n138 =  ( n30 ) ? ( LB2D_shift_x ) : ( n137 ) ;
assign n139 =  ( n23 ) ? ( n136 ) : ( n138 ) ;
assign n140 =  ( n18 ) ? ( LB2D_shift_x ) : ( n139 ) ;
assign n141 =  ( n9 ) ? ( LB2D_shift_x ) : ( n140 ) ;
assign n142 =  ( n4 ) ? ( LB2D_shift_x ) : ( n141 ) ;
assign n143 =  ( LB2D_shift_y ) < ( 10'd479 )  ;
assign n144 =  ( LB2D_shift_y ) + ( 10'd1 )  ;
assign n145 =  ( n134 ) ? ( LB2D_shift_y ) : ( n144 ) ;
assign n146 =  ( n143 ) ? ( n145 ) : ( 10'd479 ) ;
assign n147 =  ( n37 ) ? ( LB2D_shift_y ) : ( LB2D_shift_y ) ;
assign n148 =  ( n30 ) ? ( LB2D_shift_y ) : ( n147 ) ;
assign n149 =  ( n23 ) ? ( n146 ) : ( n148 ) ;
assign n150 =  ( n18 ) ? ( LB2D_shift_y ) : ( n149 ) ;
assign n151 =  ( n9 ) ? ( LB2D_shift_y ) : ( n150 ) ;
assign n152 =  ( n4 ) ? ( LB2D_shift_y ) : ( n151 ) ;
assign n153 =  ( stencil_stream_full ) == ( 1'd1 )  ;
assign n154 =  ( n153 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_0 ) ;
assign n155 = gb_fun(n154) ;
assign n156 =  ( n37 ) ? ( arg_0_TDATA ) : ( arg_0_TDATA ) ;
assign n157 =  ( n30 ) ? ( arg_0_TDATA ) : ( n156 ) ;
assign n158 =  ( n23 ) ? ( arg_0_TDATA ) : ( n157 ) ;
assign n159 =  ( n18 ) ? ( n155 ) : ( n158 ) ;
assign n160 =  ( n9 ) ? ( arg_0_TDATA ) : ( n159 ) ;
assign n161 =  ( n4 ) ? ( arg_0_TDATA ) : ( n160 ) ;
assign n162 =  ( gb_pp_it_8 ) == ( 1'd1 )  ;
assign n163 =  ( n162 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n164 =  ( n37 ) ? ( arg_0_TVALID ) : ( arg_0_TVALID ) ;
assign n165 =  ( n30 ) ? ( arg_0_TVALID ) : ( n164 ) ;
assign n166 =  ( n23 ) ? ( arg_0_TVALID ) : ( n165 ) ;
assign n167 =  ( n18 ) ? ( n163 ) : ( n166 ) ;
assign n168 =  ( n9 ) ? ( arg_0_TVALID ) : ( n167 ) ;
assign n169 =  ( n4 ) ? ( 1'd0 ) : ( n168 ) ;
assign n170 =  ( n37 ) ? ( 1'd1 ) : ( arg_1_TREADY ) ;
assign n171 =  ( n30 ) ? ( arg_1_TREADY ) : ( n170 ) ;
assign n172 =  ( n23 ) ? ( arg_1_TREADY ) : ( n171 ) ;
assign n173 =  ( n18 ) ? ( arg_1_TREADY ) : ( n172 ) ;
assign n174 =  ( n9 ) ? ( 1'd0 ) : ( n173 ) ;
assign n175 =  ( n4 ) ? ( 1'd0 ) : ( n174 ) ;
assign n176 =  ( gb_p_cnt ) + ( 19'd1 )  ;
assign n177 =  ( n176 ) == ( 19'd307200 )  ;
assign n178 =  ( n177 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n179 =  ( n37 ) ? ( gb_exit_it_1 ) : ( gb_exit_it_1 ) ;
assign n180 =  ( n30 ) ? ( gb_exit_it_1 ) : ( n179 ) ;
assign n181 =  ( n23 ) ? ( gb_exit_it_1 ) : ( n180 ) ;
assign n182 =  ( n18 ) ? ( n178 ) : ( n181 ) ;
assign n183 =  ( n9 ) ? ( gb_exit_it_1 ) : ( n182 ) ;
assign n184 =  ( n4 ) ? ( gb_exit_it_1 ) : ( n183 ) ;
assign n185 =  ( n37 ) ? ( gb_exit_it_2 ) : ( gb_exit_it_2 ) ;
assign n186 =  ( n30 ) ? ( gb_exit_it_2 ) : ( n185 ) ;
assign n187 =  ( n23 ) ? ( gb_exit_it_2 ) : ( n186 ) ;
assign n188 =  ( n18 ) ? ( gb_exit_it_1 ) : ( n187 ) ;
assign n189 =  ( n9 ) ? ( gb_exit_it_2 ) : ( n188 ) ;
assign n190 =  ( n4 ) ? ( gb_exit_it_2 ) : ( n189 ) ;
assign n191 =  ( n37 ) ? ( gb_exit_it_3 ) : ( gb_exit_it_3 ) ;
assign n192 =  ( n30 ) ? ( gb_exit_it_3 ) : ( n191 ) ;
assign n193 =  ( n23 ) ? ( gb_exit_it_3 ) : ( n192 ) ;
assign n194 =  ( n18 ) ? ( gb_exit_it_2 ) : ( n193 ) ;
assign n195 =  ( n9 ) ? ( gb_exit_it_3 ) : ( n194 ) ;
assign n196 =  ( n4 ) ? ( gb_exit_it_3 ) : ( n195 ) ;
assign n197 =  ( n37 ) ? ( gb_exit_it_4 ) : ( gb_exit_it_4 ) ;
assign n198 =  ( n30 ) ? ( gb_exit_it_4 ) : ( n197 ) ;
assign n199 =  ( n23 ) ? ( gb_exit_it_4 ) : ( n198 ) ;
assign n200 =  ( n18 ) ? ( gb_exit_it_3 ) : ( n199 ) ;
assign n201 =  ( n9 ) ? ( gb_exit_it_4 ) : ( n200 ) ;
assign n202 =  ( n4 ) ? ( gb_exit_it_4 ) : ( n201 ) ;
assign n203 =  ( n37 ) ? ( gb_exit_it_5 ) : ( gb_exit_it_5 ) ;
assign n204 =  ( n30 ) ? ( gb_exit_it_5 ) : ( n203 ) ;
assign n205 =  ( n23 ) ? ( gb_exit_it_5 ) : ( n204 ) ;
assign n206 =  ( n18 ) ? ( gb_exit_it_4 ) : ( n205 ) ;
assign n207 =  ( n9 ) ? ( gb_exit_it_5 ) : ( n206 ) ;
assign n208 =  ( n4 ) ? ( gb_exit_it_5 ) : ( n207 ) ;
assign n209 =  ( n37 ) ? ( gb_exit_it_6 ) : ( gb_exit_it_6 ) ;
assign n210 =  ( n30 ) ? ( gb_exit_it_6 ) : ( n209 ) ;
assign n211 =  ( n23 ) ? ( gb_exit_it_6 ) : ( n210 ) ;
assign n212 =  ( n18 ) ? ( gb_exit_it_5 ) : ( n211 ) ;
assign n213 =  ( n9 ) ? ( gb_exit_it_6 ) : ( n212 ) ;
assign n214 =  ( n4 ) ? ( gb_exit_it_6 ) : ( n213 ) ;
assign n215 =  ( n37 ) ? ( gb_exit_it_7 ) : ( gb_exit_it_7 ) ;
assign n216 =  ( n30 ) ? ( gb_exit_it_7 ) : ( n215 ) ;
assign n217 =  ( n23 ) ? ( gb_exit_it_7 ) : ( n216 ) ;
assign n218 =  ( n18 ) ? ( gb_exit_it_6 ) : ( n217 ) ;
assign n219 =  ( n9 ) ? ( gb_exit_it_7 ) : ( n218 ) ;
assign n220 =  ( n4 ) ? ( gb_exit_it_7 ) : ( n219 ) ;
assign n221 =  ( n37 ) ? ( gb_exit_it_8 ) : ( gb_exit_it_8 ) ;
assign n222 =  ( n30 ) ? ( gb_exit_it_8 ) : ( n221 ) ;
assign n223 =  ( n23 ) ? ( gb_exit_it_8 ) : ( n222 ) ;
assign n224 =  ( n18 ) ? ( gb_exit_it_7 ) : ( n223 ) ;
assign n225 =  ( n9 ) ? ( gb_exit_it_8 ) : ( n224 ) ;
assign n226 =  ( n4 ) ? ( gb_exit_it_8 ) : ( n225 ) ;
assign n227 =  ( gb_p_cnt ) < ( 19'd307200 )  ;
assign n228 =  ( n227 ) ? ( n176 ) : ( 19'd307200 ) ;
assign n229 =  ( n37 ) ? ( gb_p_cnt ) : ( gb_p_cnt ) ;
assign n230 =  ( n30 ) ? ( gb_p_cnt ) : ( n229 ) ;
assign n231 =  ( n23 ) ? ( gb_p_cnt ) : ( n230 ) ;
assign n232 =  ( n18 ) ? ( n228 ) : ( n231 ) ;
assign n233 =  ( n9 ) ? ( gb_p_cnt ) : ( n232 ) ;
assign n234 =  ( n4 ) ? ( gb_p_cnt ) : ( n233 ) ;
assign n235 =  ( n37 ) ? ( gb_pp_it_1 ) : ( gb_pp_it_1 ) ;
assign n236 =  ( n30 ) ? ( gb_pp_it_1 ) : ( n235 ) ;
assign n237 =  ( n23 ) ? ( gb_pp_it_1 ) : ( n236 ) ;
assign n238 =  ( n18 ) ? ( 1'd1 ) : ( n237 ) ;
assign n239 =  ( n9 ) ? ( gb_pp_it_1 ) : ( n238 ) ;
assign n240 =  ( n4 ) ? ( gb_pp_it_1 ) : ( n239 ) ;
assign n241 =  ( n37 ) ? ( gb_pp_it_2 ) : ( gb_pp_it_2 ) ;
assign n242 =  ( n30 ) ? ( gb_pp_it_2 ) : ( n241 ) ;
assign n243 =  ( n23 ) ? ( gb_pp_it_2 ) : ( n242 ) ;
assign n244 =  ( n18 ) ? ( gb_pp_it_1 ) : ( n243 ) ;
assign n245 =  ( n9 ) ? ( gb_pp_it_2 ) : ( n244 ) ;
assign n246 =  ( n4 ) ? ( gb_pp_it_2 ) : ( n245 ) ;
assign n247 =  ( n37 ) ? ( gb_pp_it_3 ) : ( gb_pp_it_3 ) ;
assign n248 =  ( n30 ) ? ( gb_pp_it_3 ) : ( n247 ) ;
assign n249 =  ( n23 ) ? ( gb_pp_it_3 ) : ( n248 ) ;
assign n250 =  ( n18 ) ? ( gb_pp_it_2 ) : ( n249 ) ;
assign n251 =  ( n9 ) ? ( gb_pp_it_3 ) : ( n250 ) ;
assign n252 =  ( n4 ) ? ( gb_pp_it_3 ) : ( n251 ) ;
assign n253 =  ( n37 ) ? ( gb_pp_it_4 ) : ( gb_pp_it_4 ) ;
assign n254 =  ( n30 ) ? ( gb_pp_it_4 ) : ( n253 ) ;
assign n255 =  ( n23 ) ? ( gb_pp_it_4 ) : ( n254 ) ;
assign n256 =  ( n18 ) ? ( gb_pp_it_3 ) : ( n255 ) ;
assign n257 =  ( n9 ) ? ( gb_pp_it_4 ) : ( n256 ) ;
assign n258 =  ( n4 ) ? ( gb_pp_it_4 ) : ( n257 ) ;
assign n259 =  ( n37 ) ? ( gb_pp_it_5 ) : ( gb_pp_it_5 ) ;
assign n260 =  ( n30 ) ? ( gb_pp_it_5 ) : ( n259 ) ;
assign n261 =  ( n23 ) ? ( gb_pp_it_5 ) : ( n260 ) ;
assign n262 =  ( n18 ) ? ( gb_pp_it_4 ) : ( n261 ) ;
assign n263 =  ( n9 ) ? ( gb_pp_it_5 ) : ( n262 ) ;
assign n264 =  ( n4 ) ? ( gb_pp_it_5 ) : ( n263 ) ;
assign n265 =  ( n37 ) ? ( gb_pp_it_6 ) : ( gb_pp_it_6 ) ;
assign n266 =  ( n30 ) ? ( gb_pp_it_6 ) : ( n265 ) ;
assign n267 =  ( n23 ) ? ( gb_pp_it_6 ) : ( n266 ) ;
assign n268 =  ( n18 ) ? ( gb_pp_it_5 ) : ( n267 ) ;
assign n269 =  ( n9 ) ? ( gb_pp_it_6 ) : ( n268 ) ;
assign n270 =  ( n4 ) ? ( gb_pp_it_6 ) : ( n269 ) ;
assign n271 =  ( n37 ) ? ( gb_pp_it_7 ) : ( gb_pp_it_7 ) ;
assign n272 =  ( n30 ) ? ( gb_pp_it_7 ) : ( n271 ) ;
assign n273 =  ( n23 ) ? ( gb_pp_it_7 ) : ( n272 ) ;
assign n274 =  ( n18 ) ? ( gb_pp_it_6 ) : ( n273 ) ;
assign n275 =  ( n9 ) ? ( gb_pp_it_7 ) : ( n274 ) ;
assign n276 =  ( n4 ) ? ( gb_pp_it_7 ) : ( n275 ) ;
assign n277 =  ( n37 ) ? ( gb_pp_it_8 ) : ( gb_pp_it_8 ) ;
assign n278 =  ( n30 ) ? ( gb_pp_it_8 ) : ( n277 ) ;
assign n279 =  ( n23 ) ? ( gb_pp_it_8 ) : ( n278 ) ;
assign n280 =  ( n18 ) ? ( gb_pp_it_7 ) : ( n279 ) ;
assign n281 =  ( n9 ) ? ( gb_pp_it_8 ) : ( n280 ) ;
assign n282 =  ( n4 ) ? ( gb_pp_it_8 ) : ( n281 ) ;
assign n283 =  ( n37 ) ? ( gb_pp_it_9 ) : ( gb_pp_it_9 ) ;
assign n284 =  ( n30 ) ? ( gb_pp_it_9 ) : ( n283 ) ;
assign n285 =  ( n23 ) ? ( gb_pp_it_9 ) : ( n284 ) ;
assign n286 =  ( n18 ) ? ( gb_pp_it_8 ) : ( n285 ) ;
assign n287 =  ( n9 ) ? ( gb_pp_it_9 ) : ( n286 ) ;
assign n288 =  ( n4 ) ? ( gb_pp_it_9 ) : ( n287 ) ;
assign n289 =  ( n37 ) ? ( LB1D_buff ) : ( in_stream_buff_0 ) ;
assign n290 =  ( n30 ) ? ( in_stream_buff_0 ) : ( n289 ) ;
assign n291 =  ( n23 ) ? ( in_stream_buff_0 ) : ( n290 ) ;
assign n292 =  ( n18 ) ? ( in_stream_buff_0 ) : ( n291 ) ;
assign n293 =  ( n9 ) ? ( in_stream_buff_0 ) : ( n292 ) ;
assign n294 =  ( n4 ) ? ( in_stream_buff_0 ) : ( n293 ) ;
assign n295 =  ( n37 ) ? ( in_stream_buff_0 ) : ( in_stream_buff_1 ) ;
assign n296 =  ( n30 ) ? ( in_stream_buff_1 ) : ( n295 ) ;
assign n297 =  ( n23 ) ? ( in_stream_buff_1 ) : ( n296 ) ;
assign n298 =  ( n18 ) ? ( in_stream_buff_1 ) : ( n297 ) ;
assign n299 =  ( n9 ) ? ( in_stream_buff_1 ) : ( n298 ) ;
assign n300 =  ( n4 ) ? ( in_stream_buff_1 ) : ( n299 ) ;
assign n301 =  ( in_stream_full ) == ( 1'd1 )  ;
assign n302 =  ( n301 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n303 =  ( n37 ) ? ( 1'd0 ) : ( in_stream_empty ) ;
assign n304 =  ( n30 ) ? ( n302 ) : ( n303 ) ;
assign n305 =  ( n23 ) ? ( in_stream_empty ) : ( n304 ) ;
assign n306 =  ( n18 ) ? ( in_stream_empty ) : ( n305 ) ;
assign n307 =  ( n9 ) ? ( in_stream_empty ) : ( n306 ) ;
assign n308 =  ( n4 ) ? ( in_stream_empty ) : ( n307 ) ;
assign n309 =  ( in_stream_empty ) == ( 1'd1 )  ;
assign n310 =  ( n309 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n311 =  ( n37 ) ? ( n310 ) : ( in_stream_full ) ;
assign n312 =  ( n30 ) ? ( 1'd0 ) : ( n311 ) ;
assign n313 =  ( n23 ) ? ( in_stream_full ) : ( n312 ) ;
assign n314 =  ( n18 ) ? ( in_stream_full ) : ( n313 ) ;
assign n315 =  ( n9 ) ? ( in_stream_full ) : ( n314 ) ;
assign n316 =  ( n4 ) ? ( in_stream_full ) : ( n315 ) ;
assign n317 =  ( n301 ) ? ( in_stream_buff_1 ) : ( in_stream_buff_0 ) ;
assign n318 =  ( LB2D_proc_w ) == ( 64'd0 )  ;
assign n319 =  (  LB2D_proc_7 [ LB2D_proc_x ] )  ;
assign n320 =  ( LB2D_proc_w ) == ( 64'd1 )  ;
assign n321 =  (  LB2D_proc_0 [ LB2D_proc_x ] )  ;
assign n322 =  ( LB2D_proc_w ) == ( 64'd2 )  ;
assign n323 =  (  LB2D_proc_1 [ LB2D_proc_x ] )  ;
assign n324 =  ( LB2D_proc_w ) == ( 64'd3 )  ;
assign n325 =  (  LB2D_proc_2 [ LB2D_proc_x ] )  ;
assign n326 =  ( LB2D_proc_w ) == ( 64'd4 )  ;
assign n327 =  (  LB2D_proc_3 [ LB2D_proc_x ] )  ;
assign n328 =  ( LB2D_proc_w ) == ( 64'd5 )  ;
assign n329 =  (  LB2D_proc_4 [ LB2D_proc_x ] )  ;
assign n330 =  ( LB2D_proc_w ) == ( 64'd6 )  ;
assign n331 =  (  LB2D_proc_5 [ LB2D_proc_x ] )  ;
assign n332 =  (  LB2D_proc_6 [ LB2D_proc_x ] )  ;
assign n333 =  ( n330 ) ? ( n331 ) : ( n332 ) ;
assign n334 =  ( n328 ) ? ( n329 ) : ( n333 ) ;
assign n335 =  ( n326 ) ? ( n327 ) : ( n334 ) ;
assign n336 =  ( n324 ) ? ( n325 ) : ( n335 ) ;
assign n337 =  ( n322 ) ? ( n323 ) : ( n336 ) ;
assign n338 =  ( n320 ) ? ( n321 ) : ( n337 ) ;
assign n339 =  ( n318 ) ? ( n319 ) : ( n338 ) ;
assign n340 =  ( n330 ) ? ( n329 ) : ( n331 ) ;
assign n341 =  ( n328 ) ? ( n327 ) : ( n340 ) ;
assign n342 =  ( n326 ) ? ( n325 ) : ( n341 ) ;
assign n343 =  ( n324 ) ? ( n323 ) : ( n342 ) ;
assign n344 =  ( n322 ) ? ( n321 ) : ( n343 ) ;
assign n345 =  ( n320 ) ? ( n319 ) : ( n344 ) ;
assign n346 =  ( n318 ) ? ( n332 ) : ( n345 ) ;
assign n347 =  ( n330 ) ? ( n327 ) : ( n329 ) ;
assign n348 =  ( n328 ) ? ( n325 ) : ( n347 ) ;
assign n349 =  ( n326 ) ? ( n323 ) : ( n348 ) ;
assign n350 =  ( n324 ) ? ( n321 ) : ( n349 ) ;
assign n351 =  ( n322 ) ? ( n319 ) : ( n350 ) ;
assign n352 =  ( n320 ) ? ( n332 ) : ( n351 ) ;
assign n353 =  ( n318 ) ? ( n331 ) : ( n352 ) ;
assign n354 =  ( n330 ) ? ( n325 ) : ( n327 ) ;
assign n355 =  ( n328 ) ? ( n323 ) : ( n354 ) ;
assign n356 =  ( n326 ) ? ( n321 ) : ( n355 ) ;
assign n357 =  ( n324 ) ? ( n319 ) : ( n356 ) ;
assign n358 =  ( n322 ) ? ( n332 ) : ( n357 ) ;
assign n359 =  ( n320 ) ? ( n331 ) : ( n358 ) ;
assign n360 =  ( n318 ) ? ( n329 ) : ( n359 ) ;
assign n361 =  ( n330 ) ? ( n323 ) : ( n325 ) ;
assign n362 =  ( n328 ) ? ( n321 ) : ( n361 ) ;
assign n363 =  ( n326 ) ? ( n319 ) : ( n362 ) ;
assign n364 =  ( n324 ) ? ( n332 ) : ( n363 ) ;
assign n365 =  ( n322 ) ? ( n331 ) : ( n364 ) ;
assign n366 =  ( n320 ) ? ( n329 ) : ( n365 ) ;
assign n367 =  ( n318 ) ? ( n327 ) : ( n366 ) ;
assign n368 =  ( n330 ) ? ( n321 ) : ( n323 ) ;
assign n369 =  ( n328 ) ? ( n319 ) : ( n368 ) ;
assign n370 =  ( n326 ) ? ( n332 ) : ( n369 ) ;
assign n371 =  ( n324 ) ? ( n331 ) : ( n370 ) ;
assign n372 =  ( n322 ) ? ( n329 ) : ( n371 ) ;
assign n373 =  ( n320 ) ? ( n327 ) : ( n372 ) ;
assign n374 =  ( n318 ) ? ( n325 ) : ( n373 ) ;
assign n375 =  ( n330 ) ? ( n319 ) : ( n321 ) ;
assign n376 =  ( n328 ) ? ( n332 ) : ( n375 ) ;
assign n377 =  ( n326 ) ? ( n331 ) : ( n376 ) ;
assign n378 =  ( n324 ) ? ( n329 ) : ( n377 ) ;
assign n379 =  ( n322 ) ? ( n327 ) : ( n378 ) ;
assign n380 =  ( n320 ) ? ( n325 ) : ( n379 ) ;
assign n381 =  ( n318 ) ? ( n323 ) : ( n380 ) ;
assign n382 =  ( n330 ) ? ( n332 ) : ( n319 ) ;
assign n383 =  ( n328 ) ? ( n331 ) : ( n382 ) ;
assign n384 =  ( n326 ) ? ( n329 ) : ( n383 ) ;
assign n385 =  ( n324 ) ? ( n327 ) : ( n384 ) ;
assign n386 =  ( n322 ) ? ( n325 ) : ( n385 ) ;
assign n387 =  ( n320 ) ? ( n323 ) : ( n386 ) ;
assign n388 =  ( n318 ) ? ( n321 ) : ( n387 ) ;
assign n389 =  { ( n381 ) , ( n388 ) }  ;
assign n390 =  { ( n374 ) , ( n389 ) }  ;
assign n391 =  { ( n367 ) , ( n390 ) }  ;
assign n392 =  { ( n360 ) , ( n391 ) }  ;
assign n393 =  { ( n353 ) , ( n392 ) }  ;
assign n394 =  { ( n346 ) , ( n393 ) }  ;
assign n395 =  { ( n339 ) , ( n394 ) }  ;
assign n396 =  { ( n317 ) , ( n395 ) }  ;
assign n397 =  ( n28 ) ? ( slice_stream_buff_0 ) : ( n396 ) ;
assign n398 =  ( n37 ) ? ( slice_stream_buff_0 ) : ( slice_stream_buff_0 ) ;
assign n399 =  ( n30 ) ? ( n397 ) : ( n398 ) ;
assign n400 =  ( n23 ) ? ( slice_stream_buff_0 ) : ( n399 ) ;
assign n401 =  ( n18 ) ? ( slice_stream_buff_0 ) : ( n400 ) ;
assign n402 =  ( n9 ) ? ( slice_stream_buff_0 ) : ( n401 ) ;
assign n403 =  ( n4 ) ? ( slice_stream_buff_0 ) : ( n402 ) ;
assign n404 =  ( n28 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n405 =  ( n37 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_1 ) ;
assign n406 =  ( n30 ) ? ( n404 ) : ( n405 ) ;
assign n407 =  ( n23 ) ? ( slice_stream_buff_1 ) : ( n406 ) ;
assign n408 =  ( n18 ) ? ( slice_stream_buff_1 ) : ( n407 ) ;
assign n409 =  ( n9 ) ? ( slice_stream_buff_1 ) : ( n408 ) ;
assign n410 =  ( n4 ) ? ( slice_stream_buff_1 ) : ( n409 ) ;
assign n411 =  ( n84 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n412 =  ( n28 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n413 =  ( n37 ) ? ( slice_stream_empty ) : ( slice_stream_empty ) ;
assign n414 =  ( n30 ) ? ( n412 ) : ( n413 ) ;
assign n415 =  ( n23 ) ? ( n411 ) : ( n414 ) ;
assign n416 =  ( n18 ) ? ( slice_stream_empty ) : ( n415 ) ;
assign n417 =  ( n9 ) ? ( slice_stream_empty ) : ( n416 ) ;
assign n418 =  ( n4 ) ? ( slice_stream_empty ) : ( n417 ) ;
assign n419 =  ( slice_stream_empty ) == ( 1'd1 )  ;
assign n420 =  ( n419 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n421 =  ( n28 ) ? ( 1'd0 ) : ( n420 ) ;
assign n422 =  ( n37 ) ? ( slice_stream_full ) : ( slice_stream_full ) ;
assign n423 =  ( n30 ) ? ( n421 ) : ( n422 ) ;
assign n424 =  ( n23 ) ? ( 1'd0 ) : ( n423 ) ;
assign n425 =  ( n18 ) ? ( slice_stream_full ) : ( n424 ) ;
assign n426 =  ( n9 ) ? ( slice_stream_full ) : ( n425 ) ;
assign n427 =  ( n4 ) ? ( slice_stream_full ) : ( n426 ) ;
assign n428 =  ( LB2D_shift_x ) >= ( 9'd8 )  ;
assign n429 = n85[71:64] ;
assign n430 = LB2D_shift_0[71:64] ;
assign n431 = LB2D_shift_1[71:64] ;
assign n432 = LB2D_shift_2[71:64] ;
assign n433 = LB2D_shift_3[71:64] ;
assign n434 = LB2D_shift_4[71:64] ;
assign n435 = LB2D_shift_5[71:64] ;
assign n436 = LB2D_shift_6[71:64] ;
assign n437 = LB2D_shift_7[71:64] ;
assign n438 =  { ( n436 ) , ( n437 ) }  ;
assign n439 =  { ( n435 ) , ( n438 ) }  ;
assign n440 =  { ( n434 ) , ( n439 ) }  ;
assign n441 =  { ( n433 ) , ( n440 ) }  ;
assign n442 =  { ( n432 ) , ( n441 ) }  ;
assign n443 =  { ( n431 ) , ( n442 ) }  ;
assign n444 =  { ( n430 ) , ( n443 ) }  ;
assign n445 =  { ( n429 ) , ( n444 ) }  ;
assign n446 = n85[63:56] ;
assign n447 = LB2D_shift_0[63:56] ;
assign n448 = LB2D_shift_1[63:56] ;
assign n449 = LB2D_shift_2[63:56] ;
assign n450 = LB2D_shift_3[63:56] ;
assign n451 = LB2D_shift_4[63:56] ;
assign n452 = LB2D_shift_5[63:56] ;
assign n453 = LB2D_shift_6[63:56] ;
assign n454 = LB2D_shift_7[63:56] ;
assign n455 =  { ( n453 ) , ( n454 ) }  ;
assign n456 =  { ( n452 ) , ( n455 ) }  ;
assign n457 =  { ( n451 ) , ( n456 ) }  ;
assign n458 =  { ( n450 ) , ( n457 ) }  ;
assign n459 =  { ( n449 ) , ( n458 ) }  ;
assign n460 =  { ( n448 ) , ( n459 ) }  ;
assign n461 =  { ( n447 ) , ( n460 ) }  ;
assign n462 =  { ( n446 ) , ( n461 ) }  ;
assign n463 = n85[55:48] ;
assign n464 = LB2D_shift_0[55:48] ;
assign n465 = LB2D_shift_1[55:48] ;
assign n466 = LB2D_shift_2[55:48] ;
assign n467 = LB2D_shift_3[55:48] ;
assign n468 = LB2D_shift_4[55:48] ;
assign n469 = LB2D_shift_5[55:48] ;
assign n470 = LB2D_shift_6[55:48] ;
assign n471 = LB2D_shift_7[55:48] ;
assign n472 =  { ( n470 ) , ( n471 ) }  ;
assign n473 =  { ( n469 ) , ( n472 ) }  ;
assign n474 =  { ( n468 ) , ( n473 ) }  ;
assign n475 =  { ( n467 ) , ( n474 ) }  ;
assign n476 =  { ( n466 ) , ( n475 ) }  ;
assign n477 =  { ( n465 ) , ( n476 ) }  ;
assign n478 =  { ( n464 ) , ( n477 ) }  ;
assign n479 =  { ( n463 ) , ( n478 ) }  ;
assign n480 = n85[47:40] ;
assign n481 = LB2D_shift_0[47:40] ;
assign n482 = LB2D_shift_1[47:40] ;
assign n483 = LB2D_shift_2[47:40] ;
assign n484 = LB2D_shift_3[47:40] ;
assign n485 = LB2D_shift_4[47:40] ;
assign n486 = LB2D_shift_5[47:40] ;
assign n487 = LB2D_shift_6[47:40] ;
assign n488 = LB2D_shift_7[47:40] ;
assign n489 =  { ( n487 ) , ( n488 ) }  ;
assign n490 =  { ( n486 ) , ( n489 ) }  ;
assign n491 =  { ( n485 ) , ( n490 ) }  ;
assign n492 =  { ( n484 ) , ( n491 ) }  ;
assign n493 =  { ( n483 ) , ( n492 ) }  ;
assign n494 =  { ( n482 ) , ( n493 ) }  ;
assign n495 =  { ( n481 ) , ( n494 ) }  ;
assign n496 =  { ( n480 ) , ( n495 ) }  ;
assign n497 = n85[39:32] ;
assign n498 = LB2D_shift_0[39:32] ;
assign n499 = LB2D_shift_1[39:32] ;
assign n500 = LB2D_shift_2[39:32] ;
assign n501 = LB2D_shift_3[39:32] ;
assign n502 = LB2D_shift_4[39:32] ;
assign n503 = LB2D_shift_5[39:32] ;
assign n504 = LB2D_shift_6[39:32] ;
assign n505 = LB2D_shift_7[39:32] ;
assign n506 =  { ( n504 ) , ( n505 ) }  ;
assign n507 =  { ( n503 ) , ( n506 ) }  ;
assign n508 =  { ( n502 ) , ( n507 ) }  ;
assign n509 =  { ( n501 ) , ( n508 ) }  ;
assign n510 =  { ( n500 ) , ( n509 ) }  ;
assign n511 =  { ( n499 ) , ( n510 ) }  ;
assign n512 =  { ( n498 ) , ( n511 ) }  ;
assign n513 =  { ( n497 ) , ( n512 ) }  ;
assign n514 = n85[31:24] ;
assign n515 = LB2D_shift_0[31:24] ;
assign n516 = LB2D_shift_1[31:24] ;
assign n517 = LB2D_shift_2[31:24] ;
assign n518 = LB2D_shift_3[31:24] ;
assign n519 = LB2D_shift_4[31:24] ;
assign n520 = LB2D_shift_5[31:24] ;
assign n521 = LB2D_shift_6[31:24] ;
assign n522 = LB2D_shift_7[31:24] ;
assign n523 =  { ( n521 ) , ( n522 ) }  ;
assign n524 =  { ( n520 ) , ( n523 ) }  ;
assign n525 =  { ( n519 ) , ( n524 ) }  ;
assign n526 =  { ( n518 ) , ( n525 ) }  ;
assign n527 =  { ( n517 ) , ( n526 ) }  ;
assign n528 =  { ( n516 ) , ( n527 ) }  ;
assign n529 =  { ( n515 ) , ( n528 ) }  ;
assign n530 =  { ( n514 ) , ( n529 ) }  ;
assign n531 = n85[23:16] ;
assign n532 = LB2D_shift_0[23:16] ;
assign n533 = LB2D_shift_1[23:16] ;
assign n534 = LB2D_shift_2[23:16] ;
assign n535 = LB2D_shift_3[23:16] ;
assign n536 = LB2D_shift_4[23:16] ;
assign n537 = LB2D_shift_5[23:16] ;
assign n538 = LB2D_shift_6[23:16] ;
assign n539 = LB2D_shift_7[23:16] ;
assign n540 =  { ( n538 ) , ( n539 ) }  ;
assign n541 =  { ( n537 ) , ( n540 ) }  ;
assign n542 =  { ( n536 ) , ( n541 ) }  ;
assign n543 =  { ( n535 ) , ( n542 ) }  ;
assign n544 =  { ( n534 ) , ( n543 ) }  ;
assign n545 =  { ( n533 ) , ( n544 ) }  ;
assign n546 =  { ( n532 ) , ( n545 ) }  ;
assign n547 =  { ( n531 ) , ( n546 ) }  ;
assign n548 = n85[15:8] ;
assign n549 = LB2D_shift_0[15:8] ;
assign n550 = LB2D_shift_1[15:8] ;
assign n551 = LB2D_shift_2[15:8] ;
assign n552 = LB2D_shift_3[15:8] ;
assign n553 = LB2D_shift_4[15:8] ;
assign n554 = LB2D_shift_5[15:8] ;
assign n555 = LB2D_shift_6[15:8] ;
assign n556 = LB2D_shift_7[15:8] ;
assign n557 =  { ( n555 ) , ( n556 ) }  ;
assign n558 =  { ( n554 ) , ( n557 ) }  ;
assign n559 =  { ( n553 ) , ( n558 ) }  ;
assign n560 =  { ( n552 ) , ( n559 ) }  ;
assign n561 =  { ( n551 ) , ( n560 ) }  ;
assign n562 =  { ( n550 ) , ( n561 ) }  ;
assign n563 =  { ( n549 ) , ( n562 ) }  ;
assign n564 =  { ( n548 ) , ( n563 ) }  ;
assign n565 = n85[7:0] ;
assign n566 = LB2D_shift_0[7:0] ;
assign n567 = LB2D_shift_1[7:0] ;
assign n568 = LB2D_shift_2[7:0] ;
assign n569 = LB2D_shift_3[7:0] ;
assign n570 = LB2D_shift_4[7:0] ;
assign n571 = LB2D_shift_5[7:0] ;
assign n572 = LB2D_shift_6[7:0] ;
assign n573 = LB2D_shift_7[7:0] ;
assign n574 =  { ( n572 ) , ( n573 ) }  ;
assign n575 =  { ( n571 ) , ( n574 ) }  ;
assign n576 =  { ( n570 ) , ( n575 ) }  ;
assign n577 =  { ( n569 ) , ( n576 ) }  ;
assign n578 =  { ( n568 ) , ( n577 ) }  ;
assign n579 =  { ( n567 ) , ( n578 ) }  ;
assign n580 =  { ( n566 ) , ( n579 ) }  ;
assign n581 =  { ( n565 ) , ( n580 ) }  ;
assign n582 =  { ( n564 ) , ( n581 ) }  ;
assign n583 =  { ( n547 ) , ( n582 ) }  ;
assign n584 =  { ( n530 ) , ( n583 ) }  ;
assign n585 =  { ( n513 ) , ( n584 ) }  ;
assign n586 =  { ( n496 ) , ( n585 ) }  ;
assign n587 =  { ( n479 ) , ( n586 ) }  ;
assign n588 =  { ( n462 ) , ( n587 ) }  ;
assign n589 =  { ( n445 ) , ( n588 ) }  ;
assign n590 =  ( n428 ) ? ( n589 ) : ( stencil_stream_buff_0 ) ;
assign n591 =  ( n37 ) ? ( stencil_stream_buff_0 ) : ( stencil_stream_buff_0 ) ;
assign n592 =  ( n30 ) ? ( stencil_stream_buff_0 ) : ( n591 ) ;
assign n593 =  ( n23 ) ? ( n590 ) : ( n592 ) ;
assign n594 =  ( n18 ) ? ( stencil_stream_buff_0 ) : ( n593 ) ;
assign n595 =  ( n9 ) ? ( stencil_stream_buff_0 ) : ( n594 ) ;
assign n596 =  ( n4 ) ? ( stencil_stream_buff_0 ) : ( n595 ) ;
assign n597 =  ( n37 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_1 ) ;
assign n598 =  ( n30 ) ? ( stencil_stream_buff_1 ) : ( n597 ) ;
assign n599 =  ( n23 ) ? ( stencil_stream_buff_0 ) : ( n598 ) ;
assign n600 =  ( n18 ) ? ( stencil_stream_buff_1 ) : ( n599 ) ;
assign n601 =  ( n9 ) ? ( stencil_stream_buff_1 ) : ( n600 ) ;
assign n602 =  ( n4 ) ? ( stencil_stream_buff_1 ) : ( n601 ) ;
assign n603 =  ( n153 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n604 =  ( n21 ) ? ( stencil_stream_empty ) : ( 1'd0 ) ;
assign n605 =  ( n37 ) ? ( stencil_stream_empty ) : ( stencil_stream_empty ) ;
assign n606 =  ( n30 ) ? ( stencil_stream_empty ) : ( n605 ) ;
assign n607 =  ( n23 ) ? ( n604 ) : ( n606 ) ;
assign n608 =  ( n18 ) ? ( n603 ) : ( n607 ) ;
assign n609 =  ( n9 ) ? ( stencil_stream_empty ) : ( n608 ) ;
assign n610 =  ( n4 ) ? ( stencil_stream_empty ) : ( n609 ) ;
assign n611 =  ( n14 ) ? ( 1'd0 ) : ( 1'd0 ) ;
assign n612 =  ( stencil_stream_empty ) == ( 1'd1 )  ;
assign n613 =  ( n612 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n614 =  ( n21 ) ? ( stencil_stream_full ) : ( n613 ) ;
assign n615 =  ( n37 ) ? ( stencil_stream_full ) : ( stencil_stream_full ) ;
assign n616 =  ( n30 ) ? ( stencil_stream_full ) : ( n615 ) ;
assign n617 =  ( n23 ) ? ( n614 ) : ( n616 ) ;
assign n618 =  ( n18 ) ? ( n611 ) : ( n617 ) ;
assign n619 =  ( n9 ) ? ( stencil_stream_full ) : ( n618 ) ;
assign n620 =  ( n4 ) ? ( stencil_stream_full ) : ( n619 ) ;
assign n621 = ~ ( n4 ) ;
assign n622 = ~ ( n9 ) ;
assign n623 =  ( n621 ) & ( n622 )  ;
assign n624 = ~ ( n18 ) ;
assign n625 =  ( n623 ) & ( n624 )  ;
assign n626 = ~ ( n23 ) ;
assign n627 =  ( n625 ) & ( n626 )  ;
assign n628 = ~ ( n30 ) ;
assign n629 =  ( n627 ) & ( n628 )  ;
assign n630 = ~ ( n37 ) ;
assign n631 =  ( n629 ) & ( n630 )  ;
assign n632 =  ( n629 ) & ( n37 )  ;
assign n633 =  ( n627 ) & ( n30 )  ;
assign n634 = ~ ( n318 ) ;
assign n635 =  ( n633 ) & ( n634 )  ;
assign n636 =  ( n633 ) & ( n318 )  ;
assign n637 =  ( n625 ) & ( n23 )  ;
assign n638 =  ( n623 ) & ( n18 )  ;
assign n639 =  ( n621 ) & ( n9 )  ;
assign LB2D_proc_0_addr0 = n636 ? (LB2D_proc_x) : (0);
assign LB2D_proc_0_data0 = n636 ? (n317) : (LB2D_proc_0[0]);
assign n640 = ~ ( n320 ) ;
assign n641 =  ( n633 ) & ( n640 )  ;
assign n642 =  ( n633 ) & ( n320 )  ;
assign LB2D_proc_1_addr0 = n642 ? (LB2D_proc_x) : (0);
assign LB2D_proc_1_data0 = n642 ? (n317) : (LB2D_proc_1[0]);
assign n643 = ~ ( n322 ) ;
assign n644 =  ( n633 ) & ( n643 )  ;
assign n645 =  ( n633 ) & ( n322 )  ;
assign LB2D_proc_2_addr0 = n645 ? (LB2D_proc_x) : (0);
assign LB2D_proc_2_data0 = n645 ? (n317) : (LB2D_proc_2[0]);
assign n646 = ~ ( n324 ) ;
assign n647 =  ( n633 ) & ( n646 )  ;
assign n648 =  ( n633 ) & ( n324 )  ;
assign LB2D_proc_3_addr0 = n648 ? (LB2D_proc_x) : (0);
assign LB2D_proc_3_data0 = n648 ? (n317) : (LB2D_proc_3[0]);
assign n649 = ~ ( n326 ) ;
assign n650 =  ( n633 ) & ( n649 )  ;
assign n651 =  ( n633 ) & ( n326 )  ;
assign LB2D_proc_4_addr0 = n651 ? (LB2D_proc_x) : (0);
assign LB2D_proc_4_data0 = n651 ? (n317) : (LB2D_proc_4[0]);
assign n652 = ~ ( n328 ) ;
assign n653 =  ( n633 ) & ( n652 )  ;
assign n654 =  ( n633 ) & ( n328 )  ;
assign LB2D_proc_5_addr0 = n654 ? (LB2D_proc_x) : (0);
assign LB2D_proc_5_data0 = n654 ? (n317) : (LB2D_proc_5[0]);
assign n655 = ~ ( n330 ) ;
assign n656 =  ( n633 ) & ( n655 )  ;
assign n657 =  ( n633 ) & ( n330 )  ;
assign LB2D_proc_6_addr0 = n657 ? (LB2D_proc_x) : (0);
assign LB2D_proc_6_data0 = n657 ? (n317) : (LB2D_proc_6[0]);
assign n658 =  ( LB2D_proc_w ) == ( 64'd7 )  ;
assign n659 = ~ ( n658 ) ;
assign n660 =  ( n633 ) & ( n659 )  ;
assign n661 =  ( n633 ) & ( n658 )  ;
assign LB2D_proc_7_addr0 = n661 ? (LB2D_proc_x) : (0);
assign LB2D_proc_7_data0 = n661 ? (n317) : (LB2D_proc_7[0]);
function [7:0] gb_fun ;
input [647:0] arg0;
    begin
//TODO: Add the specific function HERE.    end
endfunction

always @(posedge clk) begin
   if(rst) begin
       LB1D_buff <= LB1D_buff;
       LB1D_it_1 <= LB1D_it_1;
       LB1D_p_cnt <= LB1D_p_cnt;
       LB2D_proc_w <= LB2D_proc_w;
       LB2D_proc_x <= LB2D_proc_x;
       LB2D_proc_y <= LB2D_proc_y;
       LB2D_shift_0 <= LB2D_shift_0;
       LB2D_shift_1 <= LB2D_shift_1;
       LB2D_shift_2 <= LB2D_shift_2;
       LB2D_shift_3 <= LB2D_shift_3;
       LB2D_shift_4 <= LB2D_shift_4;
       LB2D_shift_5 <= LB2D_shift_5;
       LB2D_shift_6 <= LB2D_shift_6;
       LB2D_shift_7 <= LB2D_shift_7;
       LB2D_shift_x <= LB2D_shift_x;
       LB2D_shift_y <= LB2D_shift_y;
       arg_0_TDATA <= arg_0_TDATA;
       arg_0_TVALID <= arg_0_TVALID;
       arg_1_TREADY <= arg_1_TREADY;
       gb_exit_it_1 <= gb_exit_it_1;
       gb_exit_it_2 <= gb_exit_it_2;
       gb_exit_it_3 <= gb_exit_it_3;
       gb_exit_it_4 <= gb_exit_it_4;
       gb_exit_it_5 <= gb_exit_it_5;
       gb_exit_it_6 <= gb_exit_it_6;
       gb_exit_it_7 <= gb_exit_it_7;
       gb_exit_it_8 <= gb_exit_it_8;
       gb_p_cnt <= gb_p_cnt;
       gb_pp_it_1 <= gb_pp_it_1;
       gb_pp_it_2 <= gb_pp_it_2;
       gb_pp_it_3 <= gb_pp_it_3;
       gb_pp_it_4 <= gb_pp_it_4;
       gb_pp_it_5 <= gb_pp_it_5;
       gb_pp_it_6 <= gb_pp_it_6;
       gb_pp_it_7 <= gb_pp_it_7;
       gb_pp_it_8 <= gb_pp_it_8;
       gb_pp_it_9 <= gb_pp_it_9;
       in_stream_buff_0 <= in_stream_buff_0;
       in_stream_buff_1 <= in_stream_buff_1;
       in_stream_empty <= in_stream_empty;
       in_stream_full <= in_stream_full;
       slice_stream_buff_0 <= slice_stream_buff_0;
       slice_stream_buff_1 <= slice_stream_buff_1;
       slice_stream_empty <= slice_stream_empty;
       slice_stream_full <= slice_stream_full;
       stencil_stream_buff_0 <= stencil_stream_buff_0;
       stencil_stream_buff_1 <= stencil_stream_buff_1;
       stencil_stream_empty <= stencil_stream_empty;
       stencil_stream_full <= stencil_stream_full;
   end
   else if(step) begin
       LB1D_buff <= n43;
       LB1D_it_1 <= n46;
       LB1D_p_cnt <= n53;
       LB2D_proc_w <= n64;
       LB2D_proc_x <= n75;
       LB2D_proc_y <= n83;
       LB2D_shift_0 <= n91;
       LB2D_shift_1 <= n97;
       LB2D_shift_2 <= n103;
       LB2D_shift_3 <= n109;
       LB2D_shift_4 <= n115;
       LB2D_shift_5 <= n121;
       LB2D_shift_6 <= n127;
       LB2D_shift_7 <= n133;
       LB2D_shift_x <= n142;
       LB2D_shift_y <= n152;
       arg_0_TDATA <= n161;
       arg_0_TVALID <= n169;
       arg_1_TREADY <= n175;
       gb_exit_it_1 <= n184;
       gb_exit_it_2 <= n190;
       gb_exit_it_3 <= n196;
       gb_exit_it_4 <= n202;
       gb_exit_it_5 <= n208;
       gb_exit_it_6 <= n214;
       gb_exit_it_7 <= n220;
       gb_exit_it_8 <= n226;
       gb_p_cnt <= n234;
       gb_pp_it_1 <= n240;
       gb_pp_it_2 <= n246;
       gb_pp_it_3 <= n252;
       gb_pp_it_4 <= n258;
       gb_pp_it_5 <= n264;
       gb_pp_it_6 <= n270;
       gb_pp_it_7 <= n276;
       gb_pp_it_8 <= n282;
       gb_pp_it_9 <= n288;
       in_stream_buff_0 <= n294;
       in_stream_buff_1 <= n300;
       in_stream_empty <= n308;
       in_stream_full <= n316;
       slice_stream_buff_0 <= n403;
       slice_stream_buff_1 <= n410;
       slice_stream_empty <= n418;
       slice_stream_full <= n427;
       stencil_stream_buff_0 <= n596;
       stencil_stream_buff_1 <= n602;
       stencil_stream_empty <= n610;
       stencil_stream_full <= n620;
       LB2D_proc_0 [ LB2D_proc_0_addr0 ] <= LB2D_proc_0_data0;
       LB2D_proc_1 [ LB2D_proc_1_addr0 ] <= LB2D_proc_1_data0;
       LB2D_proc_2 [ LB2D_proc_2_addr0 ] <= LB2D_proc_2_data0;
       LB2D_proc_3 [ LB2D_proc_3_addr0 ] <= LB2D_proc_3_data0;
       LB2D_proc_4 [ LB2D_proc_4_addr0 ] <= LB2D_proc_4_data0;
       LB2D_proc_5 [ LB2D_proc_5_addr0 ] <= LB2D_proc_5_data0;
       LB2D_proc_6 [ LB2D_proc_6_addr0 ] <= LB2D_proc_6_data0;
       LB2D_proc_7 [ LB2D_proc_7_addr0 ] <= LB2D_proc_7_data0;
   end
end
endmodule
