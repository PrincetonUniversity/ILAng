module GB(
arg_0_TREADY,
arg_1_TDATA,
arg_1_TVALID,
LB1D_buff,
LB2D_proc_w,
LB2D_proc_x,
LB2D_proc_y,
LB2D_shift_0,
LB2D_shift_1,
LB2D_shift_2,
LB2D_shift_3,
LB2D_shift_4,
LB2D_shift_5,
LB2D_shift_6,
LB2D_shift_7,
LB2D_shift_x,
LB2D_shift_y,
arg_0_TDATA,
arg_0_TVALID,
arg_1_TREADY,
in_stream_buff_0,
in_stream_buff_1,
in_stream_empty,
in_stream_full,
slice_stream_buff_0,
slice_stream_buff_1,
slice_stream_empty,
slice_stream_full,
stencil_stream_buff_0,
stencil_stream_buff_1,
stencil_stream_empty,
stencil_stream_full,
clk,rst,
step
);
input            arg_0_TREADY;
input      [7:0] arg_1_TDATA;
input            arg_1_TVALID;
input clk;
input rst;
input step;
output      [7:0] LB1D_buff;
output     [63:0] LB2D_proc_w;
output      [8:0] LB2D_proc_x;
output      [9:0] LB2D_proc_y;
output     [71:0] LB2D_shift_0;
output     [71:0] LB2D_shift_1;
output     [71:0] LB2D_shift_2;
output     [71:0] LB2D_shift_3;
output     [71:0] LB2D_shift_4;
output     [71:0] LB2D_shift_5;
output     [71:0] LB2D_shift_6;
output     [71:0] LB2D_shift_7;
output      [8:0] LB2D_shift_x;
output      [9:0] LB2D_shift_y;
output      [7:0] arg_0_TDATA;
output            arg_0_TVALID;
output            arg_1_TREADY;
output      [7:0] in_stream_buff_0;
output      [7:0] in_stream_buff_1;
output            in_stream_empty;
output            in_stream_full;
output     [71:0] slice_stream_buff_0;
output     [71:0] slice_stream_buff_1;
output            slice_stream_empty;
output            slice_stream_full;
output    [647:0] stencil_stream_buff_0;
output    [647:0] stencil_stream_buff_1;
output            stencil_stream_empty;
output            stencil_stream_full;
reg      [7:0] LB1D_buff;
reg     [63:0] LB2D_proc_w;
reg      [8:0] LB2D_proc_x;
reg      [9:0] LB2D_proc_y;
reg     [71:0] LB2D_shift_0;
reg     [71:0] LB2D_shift_1;
reg     [71:0] LB2D_shift_2;
reg     [71:0] LB2D_shift_3;
reg     [71:0] LB2D_shift_4;
reg     [71:0] LB2D_shift_5;
reg     [71:0] LB2D_shift_6;
reg     [71:0] LB2D_shift_7;
reg      [8:0] LB2D_shift_x;
reg      [9:0] LB2D_shift_y;
reg      [7:0] arg_0_TDATA;
reg            arg_0_TVALID;
reg            arg_1_TREADY;
reg      [7:0] in_stream_buff_0;
reg      [7:0] in_stream_buff_1;
reg            in_stream_empty;
reg            in_stream_full;
reg     [71:0] slice_stream_buff_0;
reg     [71:0] slice_stream_buff_1;
reg            slice_stream_empty;
reg            slice_stream_full;
reg    [647:0] stencil_stream_buff_0;
reg    [647:0] stencil_stream_buff_1;
reg            stencil_stream_empty;
reg            stencil_stream_full;
wire            arg_0_TREADY;
wire      [7:0] arg_1_TDATA;
wire            arg_1_TVALID;
wire            n0;
wire            n1;
wire            n2;
wire            n3;
wire            n4;
wire            n5;
wire            n6;
wire            n7;
wire            n8;
wire            n9;
wire            n10;
wire            n11;
wire            n12;
wire            n13;
wire            n14;
wire            n15;
wire            n16;
wire            n17;
wire            n18;
wire            n19;
wire            n20;
wire            n21;
wire      [7:0] n22;
wire      [7:0] n23;
wire      [7:0] n24;
wire      [7:0] n25;
wire      [7:0] n26;
wire      [7:0] n27;
wire            n28;
wire            n29;
wire     [63:0] n30;
wire     [63:0] n31;
wire     [63:0] n32;
wire     [63:0] n33;
wire     [63:0] n34;
wire     [63:0] n35;
wire     [63:0] n36;
wire     [63:0] n37;
wire     [63:0] n38;
wire      [8:0] n39;
wire      [8:0] n40;
wire      [8:0] n41;
wire      [8:0] n42;
wire      [8:0] n43;
wire      [8:0] n44;
wire      [8:0] n45;
wire      [8:0] n46;
wire            n47;
wire      [9:0] n48;
wire      [9:0] n49;
wire      [9:0] n50;
wire      [9:0] n51;
wire      [9:0] n52;
wire      [9:0] n53;
wire      [9:0] n54;
wire      [9:0] n55;
wire      [9:0] n56;
wire            n57;
wire     [71:0] n58;
wire     [71:0] n59;
wire     [71:0] n60;
wire     [71:0] n61;
wire     [71:0] n62;
wire     [71:0] n63;
wire     [71:0] n64;
wire     [71:0] n65;
wire     [71:0] n66;
wire     [71:0] n67;
wire     [71:0] n68;
wire     [71:0] n69;
wire     [71:0] n70;
wire     [71:0] n71;
wire     [71:0] n72;
wire     [71:0] n73;
wire     [71:0] n74;
wire     [71:0] n75;
wire     [71:0] n76;
wire     [71:0] n77;
wire     [71:0] n78;
wire     [71:0] n79;
wire     [71:0] n80;
wire     [71:0] n81;
wire     [71:0] n82;
wire     [71:0] n83;
wire     [71:0] n84;
wire     [71:0] n85;
wire     [71:0] n86;
wire     [71:0] n87;
wire     [71:0] n88;
wire     [71:0] n89;
wire     [71:0] n90;
wire     [71:0] n91;
wire     [71:0] n92;
wire     [71:0] n93;
wire     [71:0] n94;
wire     [71:0] n95;
wire     [71:0] n96;
wire     [71:0] n97;
wire     [71:0] n98;
wire     [71:0] n99;
wire     [71:0] n100;
wire     [71:0] n101;
wire     [71:0] n102;
wire     [71:0] n103;
wire     [71:0] n104;
wire     [71:0] n105;
wire     [71:0] n106;
wire            n107;
wire      [8:0] n108;
wire      [8:0] n109;
wire      [8:0] n110;
wire      [8:0] n111;
wire      [8:0] n112;
wire      [8:0] n113;
wire      [8:0] n114;
wire      [8:0] n115;
wire      [9:0] n116;
wire      [9:0] n117;
wire      [9:0] n118;
wire      [9:0] n119;
wire      [9:0] n120;
wire      [9:0] n121;
wire            n122;
wire    [647:0] n123;
wire      [7:0] n124;
wire      [7:0] n125;
wire      [7:0] n126;
wire      [7:0] n127;
wire      [7:0] n128;
wire      [7:0] n129;
wire      [7:0] n130;
wire            n131;
wire            n132;
wire            n133;
wire            n134;
wire            n135;
wire            n136;
wire            n137;
wire            n138;
wire            n139;
wire            n140;
wire            n141;
wire            n142;
wire      [7:0] n143;
wire      [7:0] n144;
wire      [7:0] n145;
wire      [7:0] n146;
wire      [7:0] n147;
wire      [7:0] n148;
wire      [7:0] n149;
wire      [7:0] n150;
wire      [7:0] n151;
wire      [7:0] n152;
wire      [7:0] n153;
wire      [7:0] n154;
wire            n155;
wire            n156;
wire            n157;
wire            n158;
wire            n159;
wire            n160;
wire            n161;
wire            n162;
wire            n163;
wire            n164;
wire            n165;
wire            n166;
wire            n167;
wire            n168;
wire            n169;
wire            n170;
wire            n171;
wire      [7:0] n172;
wire            n173;
wire      [7:0] n174;
wire            n175;
wire      [7:0] n176;
wire            n177;
wire      [7:0] n178;
wire            n179;
wire      [7:0] n180;
wire            n181;
wire      [7:0] n182;
wire            n183;
wire      [7:0] n184;
wire            n185;
wire      [7:0] n186;
wire      [7:0] n187;
wire      [7:0] n188;
wire      [7:0] n189;
wire      [7:0] n190;
wire      [7:0] n191;
wire      [7:0] n192;
wire      [7:0] n193;
wire      [7:0] n194;
wire      [7:0] n195;
wire      [7:0] n196;
wire      [7:0] n197;
wire      [7:0] n198;
wire      [7:0] n199;
wire      [7:0] n200;
wire      [7:0] n201;
wire      [7:0] n202;
wire      [7:0] n203;
wire      [7:0] n204;
wire      [7:0] n205;
wire      [7:0] n206;
wire      [7:0] n207;
wire      [7:0] n208;
wire      [7:0] n209;
wire      [7:0] n210;
wire      [7:0] n211;
wire      [7:0] n212;
wire      [7:0] n213;
wire      [7:0] n214;
wire      [7:0] n215;
wire      [7:0] n216;
wire      [7:0] n217;
wire      [7:0] n218;
wire      [7:0] n219;
wire      [7:0] n220;
wire      [7:0] n221;
wire      [7:0] n222;
wire      [7:0] n223;
wire      [7:0] n224;
wire      [7:0] n225;
wire      [7:0] n226;
wire      [7:0] n227;
wire      [7:0] n228;
wire      [7:0] n229;
wire      [7:0] n230;
wire      [7:0] n231;
wire      [7:0] n232;
wire      [7:0] n233;
wire      [7:0] n234;
wire      [7:0] n235;
wire      [7:0] n236;
wire      [7:0] n237;
wire      [7:0] n238;
wire      [7:0] n239;
wire      [7:0] n240;
wire      [7:0] n241;
wire      [7:0] n242;
wire      [7:0] n243;
wire     [15:0] n244;
wire     [23:0] n245;
wire     [31:0] n246;
wire     [39:0] n247;
wire     [47:0] n248;
wire     [55:0] n249;
wire     [63:0] n250;
wire     [71:0] n251;
wire     [71:0] n252;
wire     [71:0] n253;
wire     [71:0] n254;
wire     [71:0] n255;
wire     [71:0] n256;
wire     [71:0] n257;
wire     [71:0] n258;
wire     [71:0] n259;
wire     [71:0] n260;
wire     [71:0] n261;
wire     [71:0] n262;
wire     [71:0] n263;
wire     [71:0] n264;
wire            n265;
wire            n266;
wire            n267;
wire            n268;
wire            n269;
wire            n270;
wire            n271;
wire            n272;
wire            n273;
wire            n274;
wire            n275;
wire            n276;
wire            n277;
wire            n278;
wire            n279;
wire            n280;
wire            n281;
wire            n282;
wire      [7:0] n283;
wire      [7:0] n284;
wire      [7:0] n285;
wire      [7:0] n286;
wire      [7:0] n287;
wire      [7:0] n288;
wire      [7:0] n289;
wire      [7:0] n290;
wire      [7:0] n291;
wire     [15:0] n292;
wire     [23:0] n293;
wire     [31:0] n294;
wire     [39:0] n295;
wire     [47:0] n296;
wire     [55:0] n297;
wire     [63:0] n298;
wire     [71:0] n299;
wire      [7:0] n300;
wire      [7:0] n301;
wire      [7:0] n302;
wire      [7:0] n303;
wire      [7:0] n304;
wire      [7:0] n305;
wire      [7:0] n306;
wire      [7:0] n307;
wire      [7:0] n308;
wire     [15:0] n309;
wire     [23:0] n310;
wire     [31:0] n311;
wire     [39:0] n312;
wire     [47:0] n313;
wire     [55:0] n314;
wire     [63:0] n315;
wire     [71:0] n316;
wire      [7:0] n317;
wire      [7:0] n318;
wire      [7:0] n319;
wire      [7:0] n320;
wire      [7:0] n321;
wire      [7:0] n322;
wire      [7:0] n323;
wire      [7:0] n324;
wire      [7:0] n325;
wire     [15:0] n326;
wire     [23:0] n327;
wire     [31:0] n328;
wire     [39:0] n329;
wire     [47:0] n330;
wire     [55:0] n331;
wire     [63:0] n332;
wire     [71:0] n333;
wire      [7:0] n334;
wire      [7:0] n335;
wire      [7:0] n336;
wire      [7:0] n337;
wire      [7:0] n338;
wire      [7:0] n339;
wire      [7:0] n340;
wire      [7:0] n341;
wire      [7:0] n342;
wire     [15:0] n343;
wire     [23:0] n344;
wire     [31:0] n345;
wire     [39:0] n346;
wire     [47:0] n347;
wire     [55:0] n348;
wire     [63:0] n349;
wire     [71:0] n350;
wire      [7:0] n351;
wire      [7:0] n352;
wire      [7:0] n353;
wire      [7:0] n354;
wire      [7:0] n355;
wire      [7:0] n356;
wire      [7:0] n357;
wire      [7:0] n358;
wire      [7:0] n359;
wire     [15:0] n360;
wire     [23:0] n361;
wire     [31:0] n362;
wire     [39:0] n363;
wire     [47:0] n364;
wire     [55:0] n365;
wire     [63:0] n366;
wire     [71:0] n367;
wire      [7:0] n368;
wire      [7:0] n369;
wire      [7:0] n370;
wire      [7:0] n371;
wire      [7:0] n372;
wire      [7:0] n373;
wire      [7:0] n374;
wire      [7:0] n375;
wire      [7:0] n376;
wire     [15:0] n377;
wire     [23:0] n378;
wire     [31:0] n379;
wire     [39:0] n380;
wire     [47:0] n381;
wire     [55:0] n382;
wire     [63:0] n383;
wire     [71:0] n384;
wire      [7:0] n385;
wire      [7:0] n386;
wire      [7:0] n387;
wire      [7:0] n388;
wire      [7:0] n389;
wire      [7:0] n390;
wire      [7:0] n391;
wire      [7:0] n392;
wire      [7:0] n393;
wire     [15:0] n394;
wire     [23:0] n395;
wire     [31:0] n396;
wire     [39:0] n397;
wire     [47:0] n398;
wire     [55:0] n399;
wire     [63:0] n400;
wire     [71:0] n401;
wire      [7:0] n402;
wire      [7:0] n403;
wire      [7:0] n404;
wire      [7:0] n405;
wire      [7:0] n406;
wire      [7:0] n407;
wire      [7:0] n408;
wire      [7:0] n409;
wire      [7:0] n410;
wire     [15:0] n411;
wire     [23:0] n412;
wire     [31:0] n413;
wire     [39:0] n414;
wire     [47:0] n415;
wire     [55:0] n416;
wire     [63:0] n417;
wire     [71:0] n418;
wire      [7:0] n419;
wire      [7:0] n420;
wire      [7:0] n421;
wire      [7:0] n422;
wire      [7:0] n423;
wire      [7:0] n424;
wire      [7:0] n425;
wire      [7:0] n426;
wire      [7:0] n427;
wire     [15:0] n428;
wire     [23:0] n429;
wire     [31:0] n430;
wire     [39:0] n431;
wire     [47:0] n432;
wire     [55:0] n433;
wire     [63:0] n434;
wire     [71:0] n435;
wire    [143:0] n436;
wire    [215:0] n437;
wire    [287:0] n438;
wire    [359:0] n439;
wire    [431:0] n440;
wire    [503:0] n441;
wire    [575:0] n442;
wire    [647:0] n443;
wire    [647:0] n444;
wire    [647:0] n445;
wire    [647:0] n446;
wire    [647:0] n447;
wire    [647:0] n448;
wire    [647:0] n449;
wire    [647:0] n450;
wire    [647:0] n451;
wire    [647:0] n452;
wire    [647:0] n453;
wire    [647:0] n454;
wire    [647:0] n455;
wire    [647:0] n456;
wire            n457;
wire            n458;
wire            n459;
wire            n460;
wire            n461;
wire            n462;
wire            n463;
wire            n464;
wire            n465;
wire            n466;
wire            n467;
wire            n468;
wire            n469;
wire            n470;
wire            n471;
wire      [8:0] LB2D_proc_0_addr0;
wire      [7:0] LB2D_proc_0_data0;
wire            n472;
wire            n473;
wire            n474;
wire            n475;
wire            n476;
wire            n477;
wire            n478;
wire            n479;
wire            n480;
wire            n481;
wire            n482;
wire            n483;
wire            n484;
wire            n485;
wire            n486;
wire            n487;
wire            n488;
wire            n489;
wire            n490;
wire      [8:0] LB2D_proc_1_addr0;
wire      [7:0] LB2D_proc_1_data0;
wire            n491;
wire            n492;
wire            n493;
wire      [8:0] LB2D_proc_2_addr0;
wire      [7:0] LB2D_proc_2_data0;
wire            n494;
wire            n495;
wire            n496;
wire      [8:0] LB2D_proc_3_addr0;
wire      [7:0] LB2D_proc_3_data0;
wire            n497;
wire            n498;
wire            n499;
wire      [8:0] LB2D_proc_4_addr0;
wire      [7:0] LB2D_proc_4_data0;
wire            n500;
wire            n501;
wire            n502;
wire      [8:0] LB2D_proc_5_addr0;
wire      [7:0] LB2D_proc_5_data0;
wire            n503;
wire            n504;
wire            n505;
wire      [8:0] LB2D_proc_6_addr0;
wire      [7:0] LB2D_proc_6_data0;
wire            n506;
wire            n507;
wire            n508;
wire      [8:0] LB2D_proc_7_addr0;
wire      [7:0] LB2D_proc_7_data0;
wire            n509;
wire            n510;
wire            n511;
wire            n512;
reg      [7:0] LB2D_proc_0[511:0];
reg      [7:0] LB2D_proc_1[511:0];
reg      [7:0] LB2D_proc_2[511:0];
reg      [7:0] LB2D_proc_3[511:0];
reg      [7:0] LB2D_proc_4[511:0];
reg      [7:0] LB2D_proc_5[511:0];
reg      [7:0] LB2D_proc_6[511:0];
reg      [7:0] LB2D_proc_7[511:0];
wire clk;
wire rst;
wire step;
assign n0 =  ( stencil_stream_empty ) == ( 1'd0 )  ;
assign n1 =  ( arg_0_TVALID ) == ( 1'd0 )  ;
assign n2 =  ( n0 ) & ( n1 )  ;
assign n3 =  ( slice_stream_empty ) == ( 1'd0 )  ;
assign n4 =  ( stencil_stream_full ) == ( 1'd0 )  ;
assign n5 =  ( n3 ) & ( n4 )  ;
assign n6 =  ( in_stream_empty ) == ( 1'd0 )  ;
assign n7 =  ( slice_stream_full ) == ( 1'd0 )  ;
assign n8 =  ( n6 ) & ( n7 )  ;
assign n9 =  ( arg_1_TREADY ) == ( 1'd0 )  ;
assign n10 =  ( in_stream_full ) == ( 1'd0 )  ;
assign n11 =  ( n9 ) & ( n10 )  ;
assign n12 =  ( arg_0_TREADY ) == ( 1'd1 )  ;
assign n13 =  ( arg_0_TVALID ) == ( 1'd1 )  ;
assign n14 =  ( n12 ) & ( n13 )  ;
assign n15 =  ( arg_1_TVALID ) == ( 1'd0 )  ;
assign n16 =  ( n14 ) & ( n15 )  ;
assign n17 =  ( arg_1_TREADY ) == ( 1'd1 )  ;
assign n18 =  ( arg_1_TVALID ) == ( 1'd1 )  ;
assign n19 =  ( n17 ) & ( n18 )  ;
assign n20 =  ( arg_0_TREADY ) == ( 1'd0 )  ;
assign n21 =  ( n19 ) & ( n20 )  ;
assign n22 =  ( n21 ) ? ( arg_1_TDATA ) : ( LB1D_buff ) ;
assign n23 =  ( n16 ) ? ( arg_1_TDATA ) : ( n22 ) ;
assign n24 =  ( n11 ) ? ( LB1D_buff ) : ( n23 ) ;
assign n25 =  ( n8 ) ? ( LB1D_buff ) : ( n24 ) ;
assign n26 =  ( n5 ) ? ( LB1D_buff ) : ( n25 ) ;
assign n27 =  ( n2 ) ? ( LB1D_buff ) : ( n26 ) ;
assign n28 =  ( LB2D_proc_w ) < ( 64'd7 )  ;
assign n29 =  ( LB2D_proc_x ) < ( 9'd487 )  ;
assign n30 =  ( LB2D_proc_w ) + ( 64'd1 )  ;
assign n31 =  ( n29 ) ? ( LB2D_proc_w ) : ( n30 ) ;
assign n32 =  ( n28 ) ? ( n31 ) : ( 64'd0 ) ;
assign n33 =  ( n21 ) ? ( LB2D_proc_w ) : ( LB2D_proc_w ) ;
assign n34 =  ( n16 ) ? ( LB2D_proc_w ) : ( n33 ) ;
assign n35 =  ( n11 ) ? ( LB2D_proc_w ) : ( n34 ) ;
assign n36 =  ( n8 ) ? ( n32 ) : ( n35 ) ;
assign n37 =  ( n5 ) ? ( LB2D_proc_w ) : ( n36 ) ;
assign n38 =  ( n2 ) ? ( LB2D_proc_w ) : ( n37 ) ;
assign n39 =  ( LB2D_proc_x ) + ( 9'd1 )  ;
assign n40 =  ( n29 ) ? ( n39 ) : ( 9'd0 ) ;
assign n41 =  ( n21 ) ? ( LB2D_proc_x ) : ( LB2D_proc_x ) ;
assign n42 =  ( n16 ) ? ( LB2D_proc_x ) : ( n41 ) ;
assign n43 =  ( n11 ) ? ( LB2D_proc_x ) : ( n42 ) ;
assign n44 =  ( n8 ) ? ( n40 ) : ( n43 ) ;
assign n45 =  ( n5 ) ? ( LB2D_proc_x ) : ( n44 ) ;
assign n46 =  ( n2 ) ? ( LB2D_proc_x ) : ( n45 ) ;
assign n47 =  ( LB2D_proc_y ) < ( 10'd487 )  ;
assign n48 =  ( LB2D_proc_y ) + ( 10'd1 )  ;
assign n49 =  ( n29 ) ? ( LB2D_proc_y ) : ( n48 ) ;
assign n50 =  ( n47 ) ? ( n49 ) : ( 10'd487 ) ;
assign n51 =  ( n21 ) ? ( LB2D_proc_y ) : ( LB2D_proc_y ) ;
assign n52 =  ( n16 ) ? ( LB2D_proc_y ) : ( n51 ) ;
assign n53 =  ( n11 ) ? ( LB2D_proc_y ) : ( n52 ) ;
assign n54 =  ( n8 ) ? ( n50 ) : ( n53 ) ;
assign n55 =  ( n5 ) ? ( LB2D_proc_y ) : ( n54 ) ;
assign n56 =  ( n2 ) ? ( LB2D_proc_y ) : ( n55 ) ;
assign n57 =  ( slice_stream_full ) == ( 1'd1 )  ;
assign n58 =  ( n57 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_0 ) ;
assign n59 =  ( n21 ) ? ( LB2D_shift_0 ) : ( LB2D_shift_0 ) ;
assign n60 =  ( n16 ) ? ( LB2D_shift_0 ) : ( n59 ) ;
assign n61 =  ( n11 ) ? ( LB2D_shift_0 ) : ( n60 ) ;
assign n62 =  ( n8 ) ? ( LB2D_shift_0 ) : ( n61 ) ;
assign n63 =  ( n5 ) ? ( n58 ) : ( n62 ) ;
assign n64 =  ( n2 ) ? ( LB2D_shift_0 ) : ( n63 ) ;
assign n65 =  ( n21 ) ? ( LB2D_shift_1 ) : ( LB2D_shift_1 ) ;
assign n66 =  ( n16 ) ? ( LB2D_shift_1 ) : ( n65 ) ;
assign n67 =  ( n11 ) ? ( LB2D_shift_1 ) : ( n66 ) ;
assign n68 =  ( n8 ) ? ( LB2D_shift_1 ) : ( n67 ) ;
assign n69 =  ( n5 ) ? ( LB2D_shift_0 ) : ( n68 ) ;
assign n70 =  ( n2 ) ? ( LB2D_shift_1 ) : ( n69 ) ;
assign n71 =  ( n21 ) ? ( LB2D_shift_2 ) : ( LB2D_shift_2 ) ;
assign n72 =  ( n16 ) ? ( LB2D_shift_2 ) : ( n71 ) ;
assign n73 =  ( n11 ) ? ( LB2D_shift_2 ) : ( n72 ) ;
assign n74 =  ( n8 ) ? ( LB2D_shift_2 ) : ( n73 ) ;
assign n75 =  ( n5 ) ? ( LB2D_shift_1 ) : ( n74 ) ;
assign n76 =  ( n2 ) ? ( LB2D_shift_2 ) : ( n75 ) ;
assign n77 =  ( n21 ) ? ( LB2D_shift_3 ) : ( LB2D_shift_3 ) ;
assign n78 =  ( n16 ) ? ( LB2D_shift_3 ) : ( n77 ) ;
assign n79 =  ( n11 ) ? ( LB2D_shift_3 ) : ( n78 ) ;
assign n80 =  ( n8 ) ? ( LB2D_shift_3 ) : ( n79 ) ;
assign n81 =  ( n5 ) ? ( LB2D_shift_2 ) : ( n80 ) ;
assign n82 =  ( n2 ) ? ( LB2D_shift_3 ) : ( n81 ) ;
assign n83 =  ( n21 ) ? ( LB2D_shift_4 ) : ( LB2D_shift_4 ) ;
assign n84 =  ( n16 ) ? ( LB2D_shift_4 ) : ( n83 ) ;
assign n85 =  ( n11 ) ? ( LB2D_shift_4 ) : ( n84 ) ;
assign n86 =  ( n8 ) ? ( LB2D_shift_4 ) : ( n85 ) ;
assign n87 =  ( n5 ) ? ( LB2D_shift_3 ) : ( n86 ) ;
assign n88 =  ( n2 ) ? ( LB2D_shift_4 ) : ( n87 ) ;
assign n89 =  ( n21 ) ? ( LB2D_shift_5 ) : ( LB2D_shift_5 ) ;
assign n90 =  ( n16 ) ? ( LB2D_shift_5 ) : ( n89 ) ;
assign n91 =  ( n11 ) ? ( LB2D_shift_5 ) : ( n90 ) ;
assign n92 =  ( n8 ) ? ( LB2D_shift_5 ) : ( n91 ) ;
assign n93 =  ( n5 ) ? ( LB2D_shift_4 ) : ( n92 ) ;
assign n94 =  ( n2 ) ? ( LB2D_shift_5 ) : ( n93 ) ;
assign n95 =  ( n21 ) ? ( LB2D_shift_6 ) : ( LB2D_shift_6 ) ;
assign n96 =  ( n16 ) ? ( LB2D_shift_6 ) : ( n95 ) ;
assign n97 =  ( n11 ) ? ( LB2D_shift_6 ) : ( n96 ) ;
assign n98 =  ( n8 ) ? ( LB2D_shift_6 ) : ( n97 ) ;
assign n99 =  ( n5 ) ? ( LB2D_shift_5 ) : ( n98 ) ;
assign n100 =  ( n2 ) ? ( LB2D_shift_6 ) : ( n99 ) ;
assign n101 =  ( n21 ) ? ( LB2D_shift_7 ) : ( LB2D_shift_7 ) ;
assign n102 =  ( n16 ) ? ( LB2D_shift_7 ) : ( n101 ) ;
assign n103 =  ( n11 ) ? ( LB2D_shift_7 ) : ( n102 ) ;
assign n104 =  ( n8 ) ? ( LB2D_shift_7 ) : ( n103 ) ;
assign n105 =  ( n5 ) ? ( LB2D_shift_6 ) : ( n104 ) ;
assign n106 =  ( n2 ) ? ( LB2D_shift_7 ) : ( n105 ) ;
assign n107 =  ( LB2D_shift_x ) < ( 9'd487 )  ;
assign n108 =  ( LB2D_shift_x ) + ( 9'd1 )  ;
assign n109 =  ( n107 ) ? ( n108 ) : ( 9'd0 ) ;
assign n110 =  ( n21 ) ? ( LB2D_shift_x ) : ( LB2D_shift_x ) ;
assign n111 =  ( n16 ) ? ( LB2D_shift_x ) : ( n110 ) ;
assign n112 =  ( n11 ) ? ( LB2D_shift_x ) : ( n111 ) ;
assign n113 =  ( n8 ) ? ( LB2D_shift_x ) : ( n112 ) ;
assign n114 =  ( n5 ) ? ( n109 ) : ( n113 ) ;
assign n115 =  ( n2 ) ? ( LB2D_shift_x ) : ( n114 ) ;
assign n116 =  ( n21 ) ? ( LB2D_shift_y ) : ( LB2D_shift_y ) ;
assign n117 =  ( n16 ) ? ( LB2D_shift_y ) : ( n116 ) ;
assign n118 =  ( n11 ) ? ( LB2D_shift_y ) : ( n117 ) ;
assign n119 =  ( n8 ) ? ( LB2D_shift_y ) : ( n118 ) ;
assign n120 =  ( n5 ) ? ( LB2D_shift_y ) : ( n119 ) ;
assign n121 =  ( n2 ) ? ( LB2D_shift_y ) : ( n120 ) ;
assign n122 =  ( stencil_stream_full ) == ( 1'd1 )  ;
assign n123 =  ( n122 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_0 ) ;
assign n124 = gb_fun(n123) ;
assign n125 =  ( n21 ) ? ( arg_0_TDATA ) : ( arg_0_TDATA ) ;
assign n126 =  ( n16 ) ? ( arg_0_TDATA ) : ( n125 ) ;
assign n127 =  ( n11 ) ? ( arg_0_TDATA ) : ( n126 ) ;
assign n128 =  ( n8 ) ? ( arg_0_TDATA ) : ( n127 ) ;
assign n129 =  ( n5 ) ? ( arg_0_TDATA ) : ( n128 ) ;
assign n130 =  ( n2 ) ? ( n124 ) : ( n129 ) ;
assign n131 =  ( n21 ) ? ( arg_0_TVALID ) : ( arg_0_TVALID ) ;
assign n132 =  ( n16 ) ? ( 1'd0 ) : ( n131 ) ;
assign n133 =  ( n11 ) ? ( arg_0_TVALID ) : ( n132 ) ;
assign n134 =  ( n8 ) ? ( arg_0_TVALID ) : ( n133 ) ;
assign n135 =  ( n5 ) ? ( arg_0_TVALID ) : ( n134 ) ;
assign n136 =  ( n2 ) ? ( 1'd1 ) : ( n135 ) ;
assign n137 =  ( n21 ) ? ( 1'd0 ) : ( arg_1_TREADY ) ;
assign n138 =  ( n16 ) ? ( 1'd0 ) : ( n137 ) ;
assign n139 =  ( n11 ) ? ( 1'd1 ) : ( n138 ) ;
assign n140 =  ( n8 ) ? ( arg_1_TREADY ) : ( n139 ) ;
assign n141 =  ( n5 ) ? ( arg_1_TREADY ) : ( n140 ) ;
assign n142 =  ( n2 ) ? ( arg_1_TREADY ) : ( n141 ) ;
assign n143 =  ( n21 ) ? ( in_stream_buff_0 ) : ( in_stream_buff_0 ) ;
assign n144 =  ( n16 ) ? ( in_stream_buff_0 ) : ( n143 ) ;
assign n145 =  ( n11 ) ? ( LB1D_buff ) : ( n144 ) ;
assign n146 =  ( n8 ) ? ( in_stream_buff_0 ) : ( n145 ) ;
assign n147 =  ( n5 ) ? ( in_stream_buff_0 ) : ( n146 ) ;
assign n148 =  ( n2 ) ? ( in_stream_buff_0 ) : ( n147 ) ;
assign n149 =  ( n21 ) ? ( in_stream_buff_1 ) : ( in_stream_buff_1 ) ;
assign n150 =  ( n16 ) ? ( in_stream_buff_1 ) : ( n149 ) ;
assign n151 =  ( n11 ) ? ( in_stream_buff_0 ) : ( n150 ) ;
assign n152 =  ( n8 ) ? ( in_stream_buff_1 ) : ( n151 ) ;
assign n153 =  ( n5 ) ? ( in_stream_buff_1 ) : ( n152 ) ;
assign n154 =  ( n2 ) ? ( in_stream_buff_1 ) : ( n153 ) ;
assign n155 =  ( in_stream_full ) == ( 1'd1 )  ;
assign n156 =  ( n155 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n157 =  ( n21 ) ? ( in_stream_empty ) : ( in_stream_empty ) ;
assign n158 =  ( n16 ) ? ( in_stream_empty ) : ( n157 ) ;
assign n159 =  ( n11 ) ? ( 1'd0 ) : ( n158 ) ;
assign n160 =  ( n8 ) ? ( n156 ) : ( n159 ) ;
assign n161 =  ( n5 ) ? ( in_stream_empty ) : ( n160 ) ;
assign n162 =  ( n2 ) ? ( in_stream_empty ) : ( n161 ) ;
assign n163 =  ( in_stream_empty ) == ( 1'd1 )  ;
assign n164 =  ( n163 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n165 =  ( n21 ) ? ( in_stream_full ) : ( in_stream_full ) ;
assign n166 =  ( n16 ) ? ( in_stream_full ) : ( n165 ) ;
assign n167 =  ( n11 ) ? ( n164 ) : ( n166 ) ;
assign n168 =  ( n8 ) ? ( 1'd0 ) : ( n167 ) ;
assign n169 =  ( n5 ) ? ( in_stream_full ) : ( n168 ) ;
assign n170 =  ( n2 ) ? ( in_stream_full ) : ( n169 ) ;
assign n171 =  ( LB2D_proc_y ) >= ( 10'd8 )  ;
assign n172 =  ( n155 ) ? ( in_stream_buff_1 ) : ( in_stream_buff_0 ) ;
assign n173 =  ( LB2D_proc_w ) == ( 64'd0 )  ;
assign n174 =  (  LB2D_proc_7 [ LB2D_proc_x ] )  ;
assign n175 =  ( LB2D_proc_w ) == ( 64'd1 )  ;
assign n176 =  (  LB2D_proc_0 [ LB2D_proc_x ] )  ;
assign n177 =  ( LB2D_proc_w ) == ( 64'd2 )  ;
assign n178 =  (  LB2D_proc_1 [ LB2D_proc_x ] )  ;
assign n179 =  ( LB2D_proc_w ) == ( 64'd3 )  ;
assign n180 =  (  LB2D_proc_2 [ LB2D_proc_x ] )  ;
assign n181 =  ( LB2D_proc_w ) == ( 64'd4 )  ;
assign n182 =  (  LB2D_proc_3 [ LB2D_proc_x ] )  ;
assign n183 =  ( LB2D_proc_w ) == ( 64'd5 )  ;
assign n184 =  (  LB2D_proc_4 [ LB2D_proc_x ] )  ;
assign n185 =  ( LB2D_proc_w ) == ( 64'd6 )  ;
assign n186 =  (  LB2D_proc_5 [ LB2D_proc_x ] )  ;
assign n187 =  (  LB2D_proc_6 [ LB2D_proc_x ] )  ;
assign n188 =  ( n185 ) ? ( n186 ) : ( n187 ) ;
assign n189 =  ( n183 ) ? ( n184 ) : ( n188 ) ;
assign n190 =  ( n181 ) ? ( n182 ) : ( n189 ) ;
assign n191 =  ( n179 ) ? ( n180 ) : ( n190 ) ;
assign n192 =  ( n177 ) ? ( n178 ) : ( n191 ) ;
assign n193 =  ( n175 ) ? ( n176 ) : ( n192 ) ;
assign n194 =  ( n173 ) ? ( n174 ) : ( n193 ) ;
assign n195 =  ( n185 ) ? ( n184 ) : ( n186 ) ;
assign n196 =  ( n183 ) ? ( n182 ) : ( n195 ) ;
assign n197 =  ( n181 ) ? ( n180 ) : ( n196 ) ;
assign n198 =  ( n179 ) ? ( n178 ) : ( n197 ) ;
assign n199 =  ( n177 ) ? ( n176 ) : ( n198 ) ;
assign n200 =  ( n175 ) ? ( n174 ) : ( n199 ) ;
assign n201 =  ( n173 ) ? ( n187 ) : ( n200 ) ;
assign n202 =  ( n185 ) ? ( n182 ) : ( n184 ) ;
assign n203 =  ( n183 ) ? ( n180 ) : ( n202 ) ;
assign n204 =  ( n181 ) ? ( n178 ) : ( n203 ) ;
assign n205 =  ( n179 ) ? ( n176 ) : ( n204 ) ;
assign n206 =  ( n177 ) ? ( n174 ) : ( n205 ) ;
assign n207 =  ( n175 ) ? ( n187 ) : ( n206 ) ;
assign n208 =  ( n173 ) ? ( n186 ) : ( n207 ) ;
assign n209 =  ( n185 ) ? ( n180 ) : ( n182 ) ;
assign n210 =  ( n183 ) ? ( n178 ) : ( n209 ) ;
assign n211 =  ( n181 ) ? ( n176 ) : ( n210 ) ;
assign n212 =  ( n179 ) ? ( n174 ) : ( n211 ) ;
assign n213 =  ( n177 ) ? ( n187 ) : ( n212 ) ;
assign n214 =  ( n175 ) ? ( n186 ) : ( n213 ) ;
assign n215 =  ( n173 ) ? ( n184 ) : ( n214 ) ;
assign n216 =  ( n185 ) ? ( n178 ) : ( n180 ) ;
assign n217 =  ( n183 ) ? ( n176 ) : ( n216 ) ;
assign n218 =  ( n181 ) ? ( n174 ) : ( n217 ) ;
assign n219 =  ( n179 ) ? ( n187 ) : ( n218 ) ;
assign n220 =  ( n177 ) ? ( n186 ) : ( n219 ) ;
assign n221 =  ( n175 ) ? ( n184 ) : ( n220 ) ;
assign n222 =  ( n173 ) ? ( n182 ) : ( n221 ) ;
assign n223 =  ( n185 ) ? ( n176 ) : ( n178 ) ;
assign n224 =  ( n183 ) ? ( n174 ) : ( n223 ) ;
assign n225 =  ( n181 ) ? ( n187 ) : ( n224 ) ;
assign n226 =  ( n179 ) ? ( n186 ) : ( n225 ) ;
assign n227 =  ( n177 ) ? ( n184 ) : ( n226 ) ;
assign n228 =  ( n175 ) ? ( n182 ) : ( n227 ) ;
assign n229 =  ( n173 ) ? ( n180 ) : ( n228 ) ;
assign n230 =  ( n185 ) ? ( n174 ) : ( n176 ) ;
assign n231 =  ( n183 ) ? ( n187 ) : ( n230 ) ;
assign n232 =  ( n181 ) ? ( n186 ) : ( n231 ) ;
assign n233 =  ( n179 ) ? ( n184 ) : ( n232 ) ;
assign n234 =  ( n177 ) ? ( n182 ) : ( n233 ) ;
assign n235 =  ( n175 ) ? ( n180 ) : ( n234 ) ;
assign n236 =  ( n173 ) ? ( n178 ) : ( n235 ) ;
assign n237 =  ( n185 ) ? ( n187 ) : ( n174 ) ;
assign n238 =  ( n183 ) ? ( n186 ) : ( n237 ) ;
assign n239 =  ( n181 ) ? ( n184 ) : ( n238 ) ;
assign n240 =  ( n179 ) ? ( n182 ) : ( n239 ) ;
assign n241 =  ( n177 ) ? ( n180 ) : ( n240 ) ;
assign n242 =  ( n175 ) ? ( n178 ) : ( n241 ) ;
assign n243 =  ( n173 ) ? ( n176 ) : ( n242 ) ;
assign n244 =  { ( n236 ) , ( n243 ) }  ;
assign n245 =  { ( n229 ) , ( n244 ) }  ;
assign n246 =  { ( n222 ) , ( n245 ) }  ;
assign n247 =  { ( n215 ) , ( n246 ) }  ;
assign n248 =  { ( n208 ) , ( n247 ) }  ;
assign n249 =  { ( n201 ) , ( n248 ) }  ;
assign n250 =  { ( n194 ) , ( n249 ) }  ;
assign n251 =  { ( n172 ) , ( n250 ) }  ;
assign n252 =  ( n171 ) ? ( n251 ) : ( slice_stream_buff_0 ) ;
assign n253 =  ( n21 ) ? ( slice_stream_buff_0 ) : ( slice_stream_buff_0 ) ;
assign n254 =  ( n16 ) ? ( slice_stream_buff_0 ) : ( n253 ) ;
assign n255 =  ( n11 ) ? ( slice_stream_buff_0 ) : ( n254 ) ;
assign n256 =  ( n8 ) ? ( n252 ) : ( n255 ) ;
assign n257 =  ( n5 ) ? ( slice_stream_buff_0 ) : ( n256 ) ;
assign n258 =  ( n2 ) ? ( slice_stream_buff_0 ) : ( n257 ) ;
assign n259 =  ( n21 ) ? ( slice_stream_buff_1 ) : ( slice_stream_buff_1 ) ;
assign n260 =  ( n16 ) ? ( slice_stream_buff_1 ) : ( n259 ) ;
assign n261 =  ( n11 ) ? ( slice_stream_buff_1 ) : ( n260 ) ;
assign n262 =  ( n8 ) ? ( slice_stream_buff_0 ) : ( n261 ) ;
assign n263 =  ( n5 ) ? ( slice_stream_buff_1 ) : ( n262 ) ;
assign n264 =  ( n2 ) ? ( slice_stream_buff_1 ) : ( n263 ) ;
assign n265 =  ( n57 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n266 =  ( n171 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n267 =  ( n21 ) ? ( slice_stream_empty ) : ( slice_stream_empty ) ;
assign n268 =  ( n16 ) ? ( slice_stream_empty ) : ( n267 ) ;
assign n269 =  ( n11 ) ? ( slice_stream_empty ) : ( n268 ) ;
assign n270 =  ( n8 ) ? ( n266 ) : ( n269 ) ;
assign n271 =  ( n5 ) ? ( n265 ) : ( n270 ) ;
assign n272 =  ( n2 ) ? ( slice_stream_empty ) : ( n271 ) ;
assign n273 =  ( slice_stream_empty ) == ( 1'd1 )  ;
assign n274 =  ( n273 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n275 =  ( n171 ) ? ( n274 ) : ( 1'd0 ) ;
assign n276 =  ( n21 ) ? ( slice_stream_full ) : ( slice_stream_full ) ;
assign n277 =  ( n16 ) ? ( slice_stream_full ) : ( n276 ) ;
assign n278 =  ( n11 ) ? ( slice_stream_full ) : ( n277 ) ;
assign n279 =  ( n8 ) ? ( n275 ) : ( n278 ) ;
assign n280 =  ( n5 ) ? ( 1'd0 ) : ( n279 ) ;
assign n281 =  ( n2 ) ? ( slice_stream_full ) : ( n280 ) ;
assign n282 =  ( LB2D_shift_x ) >= ( 9'd8 )  ;
assign n283 = n58[71:64] ;
assign n284 = LB2D_shift_0[71:64] ;
assign n285 = LB2D_shift_1[71:64] ;
assign n286 = LB2D_shift_2[71:64] ;
assign n287 = LB2D_shift_3[71:64] ;
assign n288 = LB2D_shift_4[71:64] ;
assign n289 = LB2D_shift_5[71:64] ;
assign n290 = LB2D_shift_6[71:64] ;
assign n291 = LB2D_shift_7[71:64] ;
assign n292 =  { ( n290 ) , ( n291 ) }  ;
assign n293 =  { ( n289 ) , ( n292 ) }  ;
assign n294 =  { ( n288 ) , ( n293 ) }  ;
assign n295 =  { ( n287 ) , ( n294 ) }  ;
assign n296 =  { ( n286 ) , ( n295 ) }  ;
assign n297 =  { ( n285 ) , ( n296 ) }  ;
assign n298 =  { ( n284 ) , ( n297 ) }  ;
assign n299 =  { ( n283 ) , ( n298 ) }  ;
assign n300 = n58[63:56] ;
assign n301 = LB2D_shift_0[63:56] ;
assign n302 = LB2D_shift_1[63:56] ;
assign n303 = LB2D_shift_2[63:56] ;
assign n304 = LB2D_shift_3[63:56] ;
assign n305 = LB2D_shift_4[63:56] ;
assign n306 = LB2D_shift_5[63:56] ;
assign n307 = LB2D_shift_6[63:56] ;
assign n308 = LB2D_shift_7[63:56] ;
assign n309 =  { ( n307 ) , ( n308 ) }  ;
assign n310 =  { ( n306 ) , ( n309 ) }  ;
assign n311 =  { ( n305 ) , ( n310 ) }  ;
assign n312 =  { ( n304 ) , ( n311 ) }  ;
assign n313 =  { ( n303 ) , ( n312 ) }  ;
assign n314 =  { ( n302 ) , ( n313 ) }  ;
assign n315 =  { ( n301 ) , ( n314 ) }  ;
assign n316 =  { ( n300 ) , ( n315 ) }  ;
assign n317 = n58[55:48] ;
assign n318 = LB2D_shift_0[55:48] ;
assign n319 = LB2D_shift_1[55:48] ;
assign n320 = LB2D_shift_2[55:48] ;
assign n321 = LB2D_shift_3[55:48] ;
assign n322 = LB2D_shift_4[55:48] ;
assign n323 = LB2D_shift_5[55:48] ;
assign n324 = LB2D_shift_6[55:48] ;
assign n325 = LB2D_shift_7[55:48] ;
assign n326 =  { ( n324 ) , ( n325 ) }  ;
assign n327 =  { ( n323 ) , ( n326 ) }  ;
assign n328 =  { ( n322 ) , ( n327 ) }  ;
assign n329 =  { ( n321 ) , ( n328 ) }  ;
assign n330 =  { ( n320 ) , ( n329 ) }  ;
assign n331 =  { ( n319 ) , ( n330 ) }  ;
assign n332 =  { ( n318 ) , ( n331 ) }  ;
assign n333 =  { ( n317 ) , ( n332 ) }  ;
assign n334 = n58[47:40] ;
assign n335 = LB2D_shift_0[47:40] ;
assign n336 = LB2D_shift_1[47:40] ;
assign n337 = LB2D_shift_2[47:40] ;
assign n338 = LB2D_shift_3[47:40] ;
assign n339 = LB2D_shift_4[47:40] ;
assign n340 = LB2D_shift_5[47:40] ;
assign n341 = LB2D_shift_6[47:40] ;
assign n342 = LB2D_shift_7[47:40] ;
assign n343 =  { ( n341 ) , ( n342 ) }  ;
assign n344 =  { ( n340 ) , ( n343 ) }  ;
assign n345 =  { ( n339 ) , ( n344 ) }  ;
assign n346 =  { ( n338 ) , ( n345 ) }  ;
assign n347 =  { ( n337 ) , ( n346 ) }  ;
assign n348 =  { ( n336 ) , ( n347 ) }  ;
assign n349 =  { ( n335 ) , ( n348 ) }  ;
assign n350 =  { ( n334 ) , ( n349 ) }  ;
assign n351 = n58[39:32] ;
assign n352 = LB2D_shift_0[39:32] ;
assign n353 = LB2D_shift_1[39:32] ;
assign n354 = LB2D_shift_2[39:32] ;
assign n355 = LB2D_shift_3[39:32] ;
assign n356 = LB2D_shift_4[39:32] ;
assign n357 = LB2D_shift_5[39:32] ;
assign n358 = LB2D_shift_6[39:32] ;
assign n359 = LB2D_shift_7[39:32] ;
assign n360 =  { ( n358 ) , ( n359 ) }  ;
assign n361 =  { ( n357 ) , ( n360 ) }  ;
assign n362 =  { ( n356 ) , ( n361 ) }  ;
assign n363 =  { ( n355 ) , ( n362 ) }  ;
assign n364 =  { ( n354 ) , ( n363 ) }  ;
assign n365 =  { ( n353 ) , ( n364 ) }  ;
assign n366 =  { ( n352 ) , ( n365 ) }  ;
assign n367 =  { ( n351 ) , ( n366 ) }  ;
assign n368 = n58[31:24] ;
assign n369 = LB2D_shift_0[31:24] ;
assign n370 = LB2D_shift_1[31:24] ;
assign n371 = LB2D_shift_2[31:24] ;
assign n372 = LB2D_shift_3[31:24] ;
assign n373 = LB2D_shift_4[31:24] ;
assign n374 = LB2D_shift_5[31:24] ;
assign n375 = LB2D_shift_6[31:24] ;
assign n376 = LB2D_shift_7[31:24] ;
assign n377 =  { ( n375 ) , ( n376 ) }  ;
assign n378 =  { ( n374 ) , ( n377 ) }  ;
assign n379 =  { ( n373 ) , ( n378 ) }  ;
assign n380 =  { ( n372 ) , ( n379 ) }  ;
assign n381 =  { ( n371 ) , ( n380 ) }  ;
assign n382 =  { ( n370 ) , ( n381 ) }  ;
assign n383 =  { ( n369 ) , ( n382 ) }  ;
assign n384 =  { ( n368 ) , ( n383 ) }  ;
assign n385 = n58[23:16] ;
assign n386 = LB2D_shift_0[23:16] ;
assign n387 = LB2D_shift_1[23:16] ;
assign n388 = LB2D_shift_2[23:16] ;
assign n389 = LB2D_shift_3[23:16] ;
assign n390 = LB2D_shift_4[23:16] ;
assign n391 = LB2D_shift_5[23:16] ;
assign n392 = LB2D_shift_6[23:16] ;
assign n393 = LB2D_shift_7[23:16] ;
assign n394 =  { ( n392 ) , ( n393 ) }  ;
assign n395 =  { ( n391 ) , ( n394 ) }  ;
assign n396 =  { ( n390 ) , ( n395 ) }  ;
assign n397 =  { ( n389 ) , ( n396 ) }  ;
assign n398 =  { ( n388 ) , ( n397 ) }  ;
assign n399 =  { ( n387 ) , ( n398 ) }  ;
assign n400 =  { ( n386 ) , ( n399 ) }  ;
assign n401 =  { ( n385 ) , ( n400 ) }  ;
assign n402 = n58[15:8] ;
assign n403 = LB2D_shift_0[15:8] ;
assign n404 = LB2D_shift_1[15:8] ;
assign n405 = LB2D_shift_2[15:8] ;
assign n406 = LB2D_shift_3[15:8] ;
assign n407 = LB2D_shift_4[15:8] ;
assign n408 = LB2D_shift_5[15:8] ;
assign n409 = LB2D_shift_6[15:8] ;
assign n410 = LB2D_shift_7[15:8] ;
assign n411 =  { ( n409 ) , ( n410 ) }  ;
assign n412 =  { ( n408 ) , ( n411 ) }  ;
assign n413 =  { ( n407 ) , ( n412 ) }  ;
assign n414 =  { ( n406 ) , ( n413 ) }  ;
assign n415 =  { ( n405 ) , ( n414 ) }  ;
assign n416 =  { ( n404 ) , ( n415 ) }  ;
assign n417 =  { ( n403 ) , ( n416 ) }  ;
assign n418 =  { ( n402 ) , ( n417 ) }  ;
assign n419 = n58[7:0] ;
assign n420 = LB2D_shift_0[7:0] ;
assign n421 = LB2D_shift_1[7:0] ;
assign n422 = LB2D_shift_2[7:0] ;
assign n423 = LB2D_shift_3[7:0] ;
assign n424 = LB2D_shift_4[7:0] ;
assign n425 = LB2D_shift_5[7:0] ;
assign n426 = LB2D_shift_6[7:0] ;
assign n427 = LB2D_shift_7[7:0] ;
assign n428 =  { ( n426 ) , ( n427 ) }  ;
assign n429 =  { ( n425 ) , ( n428 ) }  ;
assign n430 =  { ( n424 ) , ( n429 ) }  ;
assign n431 =  { ( n423 ) , ( n430 ) }  ;
assign n432 =  { ( n422 ) , ( n431 ) }  ;
assign n433 =  { ( n421 ) , ( n432 ) }  ;
assign n434 =  { ( n420 ) , ( n433 ) }  ;
assign n435 =  { ( n419 ) , ( n434 ) }  ;
assign n436 =  { ( n418 ) , ( n435 ) }  ;
assign n437 =  { ( n401 ) , ( n436 ) }  ;
assign n438 =  { ( n384 ) , ( n437 ) }  ;
assign n439 =  { ( n367 ) , ( n438 ) }  ;
assign n440 =  { ( n350 ) , ( n439 ) }  ;
assign n441 =  { ( n333 ) , ( n440 ) }  ;
assign n442 =  { ( n316 ) , ( n441 ) }  ;
assign n443 =  { ( n299 ) , ( n442 ) }  ;
assign n444 =  ( n282 ) ? ( n443 ) : ( stencil_stream_buff_0 ) ;
assign n445 =  ( n21 ) ? ( stencil_stream_buff_0 ) : ( stencil_stream_buff_0 ) ;
assign n446 =  ( n16 ) ? ( stencil_stream_buff_0 ) : ( n445 ) ;
assign n447 =  ( n11 ) ? ( stencil_stream_buff_0 ) : ( n446 ) ;
assign n448 =  ( n8 ) ? ( stencil_stream_buff_0 ) : ( n447 ) ;
assign n449 =  ( n5 ) ? ( n444 ) : ( n448 ) ;
assign n450 =  ( n2 ) ? ( stencil_stream_buff_0 ) : ( n449 ) ;
assign n451 =  ( n21 ) ? ( stencil_stream_buff_1 ) : ( stencil_stream_buff_1 ) ;
assign n452 =  ( n16 ) ? ( stencil_stream_buff_1 ) : ( n451 ) ;
assign n453 =  ( n11 ) ? ( stencil_stream_buff_1 ) : ( n452 ) ;
assign n454 =  ( n8 ) ? ( stencil_stream_buff_1 ) : ( n453 ) ;
assign n455 =  ( n5 ) ? ( stencil_stream_buff_0 ) : ( n454 ) ;
assign n456 =  ( n2 ) ? ( stencil_stream_buff_1 ) : ( n455 ) ;
assign n457 =  ( n122 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n458 =  ( n21 ) ? ( stencil_stream_empty ) : ( stencil_stream_empty ) ;
assign n459 =  ( n16 ) ? ( stencil_stream_empty ) : ( n458 ) ;
assign n460 =  ( n11 ) ? ( stencil_stream_empty ) : ( n459 ) ;
assign n461 =  ( n8 ) ? ( stencil_stream_empty ) : ( n460 ) ;
assign n462 =  ( n2 ) ? ( n457 ) : ( n461 ) ;
assign n463 =  ( stencil_stream_empty ) == ( 1'd1 )  ;
assign n464 =  ( n463 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n465 =  ( n282 ) ? ( n464 ) : ( 1'd0 ) ;
assign n466 =  ( n21 ) ? ( stencil_stream_full ) : ( stencil_stream_full ) ;
assign n467 =  ( n16 ) ? ( stencil_stream_full ) : ( n466 ) ;
assign n468 =  ( n11 ) ? ( stencil_stream_full ) : ( n467 ) ;
assign n469 =  ( n8 ) ? ( stencil_stream_full ) : ( n468 ) ;
assign n470 =  ( n5 ) ? ( n465 ) : ( n469 ) ;
assign n471 =  ( n2 ) ? ( 1'd0 ) : ( n470 ) ;
assign n472 = ~ ( n2 ) ;
assign n473 = ~ ( n5 ) ;
assign n474 =  ( n472 ) & ( n473 )  ;
assign n475 = ~ ( n8 ) ;
assign n476 =  ( n474 ) & ( n475 )  ;
assign n477 = ~ ( n11 ) ;
assign n478 =  ( n476 ) & ( n477 )  ;
assign n479 = ~ ( n16 ) ;
assign n480 =  ( n478 ) & ( n479 )  ;
assign n481 = ~ ( n21 ) ;
assign n482 =  ( n480 ) & ( n481 )  ;
assign n483 =  ( n480 ) & ( n21 )  ;
assign n484 =  ( n478 ) & ( n16 )  ;
assign n485 =  ( n476 ) & ( n11 )  ;
assign n486 =  ( n474 ) & ( n8 )  ;
assign n487 = ~ ( n173 ) ;
assign n488 =  ( n486 ) & ( n487 )  ;
assign n489 =  ( n486 ) & ( n173 )  ;
assign n490 =  ( n472 ) & ( n5 )  ;
assign LB2D_proc_0_addr0 = n489 ? (LB2D_proc_x) : (0);
assign LB2D_proc_0_data0 = n489 ? (n172) : (LB2D_proc_0[0]);
assign n491 = ~ ( n175 ) ;
assign n492 =  ( n486 ) & ( n491 )  ;
assign n493 =  ( n486 ) & ( n175 )  ;
assign LB2D_proc_1_addr0 = n493 ? (LB2D_proc_x) : (0);
assign LB2D_proc_1_data0 = n493 ? (n172) : (LB2D_proc_1[0]);
assign n494 = ~ ( n177 ) ;
assign n495 =  ( n486 ) & ( n494 )  ;
assign n496 =  ( n486 ) & ( n177 )  ;
assign LB2D_proc_2_addr0 = n496 ? (LB2D_proc_x) : (0);
assign LB2D_proc_2_data0 = n496 ? (n172) : (LB2D_proc_2[0]);
assign n497 = ~ ( n179 ) ;
assign n498 =  ( n486 ) & ( n497 )  ;
assign n499 =  ( n486 ) & ( n179 )  ;
assign LB2D_proc_3_addr0 = n499 ? (LB2D_proc_x) : (0);
assign LB2D_proc_3_data0 = n499 ? (n172) : (LB2D_proc_3[0]);
assign n500 = ~ ( n181 ) ;
assign n501 =  ( n486 ) & ( n500 )  ;
assign n502 =  ( n486 ) & ( n181 )  ;
assign LB2D_proc_4_addr0 = n502 ? (LB2D_proc_x) : (0);
assign LB2D_proc_4_data0 = n502 ? (n172) : (LB2D_proc_4[0]);
assign n503 = ~ ( n183 ) ;
assign n504 =  ( n486 ) & ( n503 )  ;
assign n505 =  ( n486 ) & ( n183 )  ;
assign LB2D_proc_5_addr0 = n505 ? (LB2D_proc_x) : (0);
assign LB2D_proc_5_data0 = n505 ? (n172) : (LB2D_proc_5[0]);
assign n506 = ~ ( n185 ) ;
assign n507 =  ( n486 ) & ( n506 )  ;
assign n508 =  ( n486 ) & ( n185 )  ;
assign LB2D_proc_6_addr0 = n508 ? (LB2D_proc_x) : (0);
assign LB2D_proc_6_data0 = n508 ? (n172) : (LB2D_proc_6[0]);
assign n509 =  ( LB2D_proc_w ) == ( 64'd7 )  ;
assign n510 = ~ ( n509 ) ;
assign n511 =  ( n486 ) & ( n510 )  ;
assign n512 =  ( n486 ) & ( n509 )  ;
assign LB2D_proc_7_addr0 = n512 ? (LB2D_proc_x) : (0);
assign LB2D_proc_7_data0 = n512 ? (n172) : (LB2D_proc_7[0]);
function [7:0] gb_fun ;
input [647:0] arg0;
    begin
//TODO: Add the specific function HERE.    end
endfunction

always @(posedge clk) begin
   if(rst) begin
       LB1D_buff <= LB1D_buff;
       LB2D_proc_w <= LB2D_proc_w;
       LB2D_proc_x <= LB2D_proc_x;
       LB2D_proc_y <= LB2D_proc_y;
       LB2D_shift_0 <= LB2D_shift_0;
       LB2D_shift_1 <= LB2D_shift_1;
       LB2D_shift_2 <= LB2D_shift_2;
       LB2D_shift_3 <= LB2D_shift_3;
       LB2D_shift_4 <= LB2D_shift_4;
       LB2D_shift_5 <= LB2D_shift_5;
       LB2D_shift_6 <= LB2D_shift_6;
       LB2D_shift_7 <= LB2D_shift_7;
       LB2D_shift_x <= LB2D_shift_x;
       LB2D_shift_y <= LB2D_shift_y;
       arg_0_TDATA <= arg_0_TDATA;
       arg_0_TVALID <= arg_0_TVALID;
       arg_1_TREADY <= arg_1_TREADY;
       in_stream_buff_0 <= in_stream_buff_0;
       in_stream_buff_1 <= in_stream_buff_1;
       in_stream_empty <= in_stream_empty;
       in_stream_full <= in_stream_full;
       slice_stream_buff_0 <= slice_stream_buff_0;
       slice_stream_buff_1 <= slice_stream_buff_1;
       slice_stream_empty <= slice_stream_empty;
       slice_stream_full <= slice_stream_full;
       stencil_stream_buff_0 <= stencil_stream_buff_0;
       stencil_stream_buff_1 <= stencil_stream_buff_1;
       stencil_stream_empty <= stencil_stream_empty;
       stencil_stream_full <= stencil_stream_full;
   end
   else if(step) begin
       LB1D_buff <= n27;
       LB2D_proc_w <= n38;
       LB2D_proc_x <= n46;
       LB2D_proc_y <= n56;
       LB2D_shift_0 <= n64;
       LB2D_shift_1 <= n70;
       LB2D_shift_2 <= n76;
       LB2D_shift_3 <= n82;
       LB2D_shift_4 <= n88;
       LB2D_shift_5 <= n94;
       LB2D_shift_6 <= n100;
       LB2D_shift_7 <= n106;
       LB2D_shift_x <= n115;
       LB2D_shift_y <= n121;
       arg_0_TDATA <= n130;
       arg_0_TVALID <= n136;
       arg_1_TREADY <= n142;
       in_stream_buff_0 <= n148;
       in_stream_buff_1 <= n154;
       in_stream_empty <= n162;
       in_stream_full <= n170;
       slice_stream_buff_0 <= n258;
       slice_stream_buff_1 <= n264;
       slice_stream_empty <= n272;
       slice_stream_full <= n281;
       stencil_stream_buff_0 <= n450;
       stencil_stream_buff_1 <= n456;
       stencil_stream_empty <= n462;
       stencil_stream_full <= n471;
       LB2D_proc_0 [ LB2D_proc_0_addr0 ] <= LB2D_proc_0_data0;
       LB2D_proc_1 [ LB2D_proc_1_addr0 ] <= LB2D_proc_1_data0;
       LB2D_proc_2 [ LB2D_proc_2_addr0 ] <= LB2D_proc_2_data0;
       LB2D_proc_3 [ LB2D_proc_3_addr0 ] <= LB2D_proc_3_data0;
       LB2D_proc_4 [ LB2D_proc_4_addr0 ] <= LB2D_proc_4_data0;
       LB2D_proc_5 [ LB2D_proc_5_addr0 ] <= LB2D_proc_5_data0;
       LB2D_proc_6 [ LB2D_proc_6_addr0 ] <= LB2D_proc_6_data0;
       LB2D_proc_7 [ LB2D_proc_7_addr0 ] <= LB2D_proc_7_data0;
   end
end
endmodule
