module GB(
arg_0_TREADY,
arg_1_TDATA,
arg_1_TVALID,
RAM_w,
RAM_x,
RAM_y,
arg_0_TDATA,
arg_0_TVALID,
arg_1_TREADY,
cur_pix,
pre_pix,
proc_in,
st_ready,
stencil_0,
stencil_1,
stencil_2,
stencil_3,
stencil_4,
stencil_5,
stencil_6,
stencil_7,
stencil_8,
clk,rst,
step
);
input            arg_0_TREADY;
input      [7:0] arg_1_TDATA;
input            arg_1_TVALID;
input clk;
input rst;
input step;
output      [2:0] RAM_w;
output      [8:0] RAM_x;
output      [9:0] RAM_y;
output      [7:0] arg_0_TDATA;
output            arg_0_TVALID;
output            arg_1_TREADY;
output      [7:0] cur_pix;
output      [7:0] pre_pix;
output    [647:0] proc_in;
output            st_ready;
output     [71:0] stencil_0;
output     [71:0] stencil_1;
output     [71:0] stencil_2;
output     [71:0] stencil_3;
output     [71:0] stencil_4;
output     [71:0] stencil_5;
output     [71:0] stencil_6;
output     [71:0] stencil_7;
output     [71:0] stencil_8;
reg      [2:0] RAM_w;
reg      [8:0] RAM_x;
reg      [9:0] RAM_y;
reg      [7:0] arg_0_TDATA;
reg            arg_0_TVALID;
reg            arg_1_TREADY;
reg      [7:0] cur_pix;
reg      [7:0] pre_pix;
reg    [647:0] proc_in;
reg            st_ready;
reg     [71:0] stencil_0;
reg     [71:0] stencil_1;
reg     [71:0] stencil_2;
reg     [71:0] stencil_3;
reg     [71:0] stencil_4;
reg     [71:0] stencil_5;
reg     [71:0] stencil_6;
reg     [71:0] stencil_7;
reg     [71:0] stencil_8;
wire            arg_0_TREADY;
wire      [7:0] arg_1_TDATA;
wire            arg_1_TVALID;
wire            n0;
wire            n1;
wire            n2;
wire            n3;
wire            n4;
wire            n5;
wire            n6;
wire            n7;
wire            n8;
wire            n9;
wire            n10;
wire            n11;
wire            n12;
wire            n13;
wire            n14;
wire            n15;
wire            n16;
wire            n17;
wire      [2:0] n18;
wire      [2:0] n19;
wire      [2:0] n20;
wire            n21;
wire            n22;
wire            n23;
wire            n24;
wire            n25;
wire      [2:0] n26;
wire      [2:0] n27;
wire      [2:0] n28;
wire      [2:0] n29;
wire      [8:0] n30;
wire      [8:0] n31;
wire      [8:0] n32;
wire      [8:0] n33;
wire      [8:0] n34;
wire      [8:0] n35;
wire            n36;
wire      [9:0] n37;
wire      [9:0] n38;
wire      [9:0] n39;
wire      [9:0] n40;
wire      [9:0] n41;
wire      [9:0] n42;
wire      [9:0] n43;
wire            n44;
wire      [7:0] n45;
wire      [7:0] n46;
wire      [7:0] n47;
wire      [7:0] n48;
wire      [7:0] n49;
wire      [7:0] n50;
wire      [7:0] n51;
wire      [7:0] n52;
wire      [7:0] n53;
wire     [15:0] n54;
wire     [23:0] n55;
wire     [31:0] n56;
wire     [39:0] n57;
wire     [47:0] n58;
wire     [55:0] n59;
wire     [63:0] n60;
wire     [71:0] n61;
wire      [7:0] n62;
wire      [7:0] n63;
wire      [7:0] n64;
wire      [7:0] n65;
wire      [7:0] n66;
wire      [7:0] n67;
wire      [7:0] n68;
wire      [7:0] n69;
wire      [7:0] n70;
wire     [15:0] n71;
wire     [23:0] n72;
wire     [31:0] n73;
wire     [39:0] n74;
wire     [47:0] n75;
wire     [55:0] n76;
wire     [63:0] n77;
wire     [71:0] n78;
wire      [7:0] n79;
wire      [7:0] n80;
wire      [7:0] n81;
wire      [7:0] n82;
wire      [7:0] n83;
wire      [7:0] n84;
wire      [7:0] n85;
wire      [7:0] n86;
wire      [7:0] n87;
wire     [15:0] n88;
wire     [23:0] n89;
wire     [31:0] n90;
wire     [39:0] n91;
wire     [47:0] n92;
wire     [55:0] n93;
wire     [63:0] n94;
wire     [71:0] n95;
wire      [7:0] n96;
wire      [7:0] n97;
wire      [7:0] n98;
wire      [7:0] n99;
wire      [7:0] n100;
wire      [7:0] n101;
wire      [7:0] n102;
wire      [7:0] n103;
wire      [7:0] n104;
wire     [15:0] n105;
wire     [23:0] n106;
wire     [31:0] n107;
wire     [39:0] n108;
wire     [47:0] n109;
wire     [55:0] n110;
wire     [63:0] n111;
wire     [71:0] n112;
wire      [7:0] n113;
wire      [7:0] n114;
wire      [7:0] n115;
wire      [7:0] n116;
wire      [7:0] n117;
wire      [7:0] n118;
wire      [7:0] n119;
wire      [7:0] n120;
wire      [7:0] n121;
wire     [15:0] n122;
wire     [23:0] n123;
wire     [31:0] n124;
wire     [39:0] n125;
wire     [47:0] n126;
wire     [55:0] n127;
wire     [63:0] n128;
wire     [71:0] n129;
wire      [7:0] n130;
wire      [7:0] n131;
wire      [7:0] n132;
wire      [7:0] n133;
wire      [7:0] n134;
wire      [7:0] n135;
wire      [7:0] n136;
wire      [7:0] n137;
wire      [7:0] n138;
wire     [15:0] n139;
wire     [23:0] n140;
wire     [31:0] n141;
wire     [39:0] n142;
wire     [47:0] n143;
wire     [55:0] n144;
wire     [63:0] n145;
wire     [71:0] n146;
wire      [7:0] n147;
wire      [7:0] n148;
wire      [7:0] n149;
wire      [7:0] n150;
wire      [7:0] n151;
wire      [7:0] n152;
wire      [7:0] n153;
wire      [7:0] n154;
wire      [7:0] n155;
wire     [15:0] n156;
wire     [23:0] n157;
wire     [31:0] n158;
wire     [39:0] n159;
wire     [47:0] n160;
wire     [55:0] n161;
wire     [63:0] n162;
wire     [71:0] n163;
wire      [7:0] n164;
wire      [7:0] n165;
wire      [7:0] n166;
wire      [7:0] n167;
wire      [7:0] n168;
wire      [7:0] n169;
wire      [7:0] n170;
wire      [7:0] n171;
wire      [7:0] n172;
wire     [15:0] n173;
wire     [23:0] n174;
wire     [31:0] n175;
wire     [39:0] n176;
wire     [47:0] n177;
wire     [55:0] n178;
wire     [63:0] n179;
wire     [71:0] n180;
wire      [7:0] n181;
wire      [7:0] n182;
wire      [7:0] n183;
wire      [7:0] n184;
wire      [7:0] n185;
wire      [7:0] n186;
wire      [7:0] n187;
wire      [7:0] n188;
wire      [7:0] n189;
wire     [15:0] n190;
wire     [23:0] n191;
wire     [31:0] n192;
wire     [39:0] n193;
wire     [47:0] n194;
wire     [55:0] n195;
wire     [63:0] n196;
wire     [71:0] n197;
wire    [143:0] n198;
wire    [215:0] n199;
wire    [287:0] n200;
wire    [359:0] n201;
wire    [431:0] n202;
wire    [503:0] n203;
wire    [575:0] n204;
wire    [647:0] n205;
wire    [647:0] n206;
wire      [7:0] n207;
wire      [7:0] n208;
wire      [7:0] n209;
wire      [7:0] n210;
wire      [7:0] n211;
wire            n212;
wire            n213;
wire            n214;
wire            n215;
wire            n216;
wire            n217;
wire            n218;
wire            n219;
wire            n220;
wire            n221;
wire            n222;
wire            n223;
wire      [9:0] n224;
wire            n225;
wire            n226;
wire            n227;
wire            n228;
wire            n229;
wire            n230;
wire            n231;
wire            n232;
wire      [7:0] n233;
wire      [7:0] n234;
wire      [7:0] n235;
wire      [7:0] n236;
wire      [7:0] n237;
wire      [7:0] n238;
wire      [7:0] n239;
wire    [647:0] n240;
wire    [647:0] n241;
wire    [647:0] n242;
wire            n243;
wire            n244;
wire            n245;
wire            n246;
wire     [71:0] n247;
wire     [71:0] n248;
wire     [71:0] n249;
wire     [71:0] n250;
wire     [71:0] n251;
wire     [71:0] n252;
wire     [71:0] n253;
wire     [71:0] n254;
wire     [71:0] n255;
wire     [71:0] n256;
wire     [71:0] n257;
wire     [71:0] n258;
wire     [71:0] n259;
wire     [71:0] n260;
wire     [71:0] n261;
wire     [71:0] n262;
wire     [71:0] n263;
wire     [71:0] n264;
wire     [71:0] n265;
wire     [71:0] n266;
wire     [71:0] n267;
wire     [71:0] n268;
wire     [71:0] n269;
wire     [71:0] n270;
wire     [71:0] n271;
wire     [71:0] n272;
wire     [71:0] n273;
wire     [71:0] n274;
wire     [71:0] n275;
wire     [71:0] n276;
wire     [71:0] n277;
wire     [71:0] n278;
wire     [71:0] n279;
wire     [71:0] n280;
wire     [71:0] n281;
wire     [71:0] n282;
wire     [71:0] n283;
wire     [71:0] n284;
wire     [71:0] n285;
wire     [71:0] n286;
wire            n287;
wire      [8:0] n288;
wire      [7:0] n289;
wire            n290;
wire            n291;
wire            n292;
wire            n293;
wire            n294;
wire            n295;
wire      [7:0] n296;
wire      [7:0] n297;
wire      [7:0] n298;
wire      [7:0] n299;
wire      [7:0] n300;
wire      [7:0] n301;
wire      [7:0] n302;
wire      [7:0] n303;
wire      [7:0] n304;
wire      [7:0] n305;
wire      [7:0] n306;
wire      [7:0] n307;
wire      [7:0] n308;
wire      [7:0] n309;
wire      [7:0] n310;
wire      [7:0] n311;
wire      [7:0] n312;
wire      [7:0] n313;
wire      [7:0] n314;
wire      [7:0] n315;
wire      [7:0] n316;
wire      [7:0] n317;
wire      [7:0] n318;
wire      [7:0] n319;
wire      [7:0] n320;
wire      [7:0] n321;
wire      [7:0] n322;
wire      [7:0] n323;
wire      [7:0] n324;
wire      [7:0] n325;
wire      [7:0] n326;
wire      [7:0] n327;
wire      [7:0] n328;
wire      [7:0] n329;
wire      [7:0] n330;
wire      [7:0] n331;
wire      [7:0] n332;
wire      [7:0] n333;
wire      [7:0] n334;
wire      [7:0] n335;
wire      [7:0] n336;
wire      [7:0] n337;
wire      [7:0] n338;
wire      [7:0] n339;
wire      [7:0] n340;
wire      [7:0] n341;
wire      [7:0] n342;
wire      [7:0] n343;
wire      [7:0] n344;
wire      [7:0] n345;
wire      [7:0] n346;
wire      [7:0] n347;
wire      [7:0] n348;
wire      [7:0] n349;
wire      [7:0] n350;
wire      [7:0] n351;
wire      [7:0] n352;
wire      [7:0] n353;
wire      [7:0] n354;
wire      [7:0] n355;
wire      [7:0] n356;
wire      [7:0] n357;
wire      [7:0] n358;
wire     [15:0] n359;
wire     [23:0] n360;
wire     [31:0] n361;
wire     [39:0] n362;
wire     [47:0] n363;
wire     [55:0] n364;
wire     [63:0] n365;
wire     [71:0] n366;
wire     [71:0] n367;
wire     [71:0] n368;
wire     [71:0] n369;
wire     [71:0] n370;
wire     [71:0] n371;
wire      [8:0] RAM_0_addr0;
wire      [7:0] RAM_0_data0;
wire            n372;
wire            n373;
wire            n374;
wire            n375;
wire            n376;
wire            n377;
wire            n378;
wire            n379;
wire            n380;
wire            n381;
wire            n382;
wire            n383;
wire            n384;
wire      [8:0] RAM_1_addr0;
wire      [7:0] RAM_1_data0;
wire            n385;
wire            n386;
wire            n387;
wire      [8:0] RAM_2_addr0;
wire      [7:0] RAM_2_data0;
wire            n388;
wire            n389;
wire            n390;
wire      [8:0] RAM_3_addr0;
wire      [7:0] RAM_3_data0;
wire            n391;
wire            n392;
wire            n393;
wire      [8:0] RAM_4_addr0;
wire      [7:0] RAM_4_data0;
wire            n394;
wire            n395;
wire            n396;
wire      [8:0] RAM_5_addr0;
wire      [7:0] RAM_5_data0;
wire            n397;
wire            n398;
wire            n399;
wire      [8:0] RAM_6_addr0;
wire      [7:0] RAM_6_data0;
wire            n400;
wire            n401;
wire            n402;
wire      [8:0] RAM_7_addr0;
wire      [7:0] RAM_7_data0;
wire            n403;
wire            n404;
wire            n405;
reg      [7:0] RAM_0[511:0];
reg      [7:0] RAM_1[511:0];
reg      [7:0] RAM_2[511:0];
reg      [7:0] RAM_3[511:0];
reg      [7:0] RAM_4[511:0];
reg      [7:0] RAM_5[511:0];
reg      [7:0] RAM_6[511:0];
reg      [7:0] RAM_7[511:0];
wire clk;
wire rst;
wire step;
assign n0 =  ( arg_1_TREADY ) == ( 1'd0 )  ;
assign n1 =  ( arg_0_TVALID ) == ( 1'd0 )  ;
assign n2 =  ( n0 ) & ( n1 )  ;
assign n3 =  ( arg_0_TREADY ) == ( 1'd0 )  ;
assign n4 =  ( n2 ) & ( n3 )  ;
assign n5 =  ( st_ready ) == ( 1'd0 )  ;
assign n6 =  ( n4 ) & ( n5 )  ;
assign n7 =  ( st_ready ) == ( 1'd1 )  ;
assign n8 =  ( n4 ) & ( n7 )  ;
assign n9 =  ( RAM_x ) == ( 9'd0 )  ;
assign n10 =  ( n8 ) & ( n9 )  ;
assign n11 =  ( RAM_y ) == ( 10'd0 )  ;
assign n12 =  ( n10 ) & ( n11 )  ;
assign n13 =  ( n9 ) & ( n11 )  ;
assign n14 = ~ ( n13 ) ;
assign n15 =  ( n8 ) & ( n14 )  ;
assign n16 =  ( RAM_x ) == ( 9'd488 )  ;
assign n17 =  ( RAM_w ) == ( 3'd7 )  ;
assign n18 =  ( RAM_w ) + ( 3'd1 )  ;
assign n19 =  ( n17 ) ? ( 3'd0 ) : ( n18 ) ;
assign n20 =  ( n16 ) ? ( n19 ) : ( RAM_w ) ;
assign n21 =  ( arg_1_TVALID ) == ( 1'd1 )  ;
assign n22 =  ( arg_1_TREADY ) == ( 1'd1 )  ;
assign n23 =  ( n21 ) & ( n22 )  ;
assign n24 =  ( n23 ) & ( n1 )  ;
assign n25 =  ( n24 ) & ( n3 )  ;
assign n26 =  ( n25 ) ? ( RAM_w ) : ( RAM_w ) ;
assign n27 =  ( n15 ) ? ( n20 ) : ( n26 ) ;
assign n28 =  ( n12 ) ? ( RAM_w ) : ( n27 ) ;
assign n29 =  ( n6 ) ? ( RAM_w ) : ( n28 ) ;
assign n30 =  ( RAM_x ) + ( 9'd1 )  ;
assign n31 =  ( n16 ) ? ( 9'd1 ) : ( n30 ) ;
assign n32 =  ( n25 ) ? ( RAM_x ) : ( RAM_x ) ;
assign n33 =  ( n15 ) ? ( n31 ) : ( n32 ) ;
assign n34 =  ( n12 ) ? ( 9'd1 ) : ( n33 ) ;
assign n35 =  ( n6 ) ? ( RAM_x ) : ( n34 ) ;
assign n36 =  ( RAM_y ) == ( 10'd648 )  ;
assign n37 =  ( RAM_y ) + ( 10'd1 )  ;
assign n38 =  ( n36 ) ? ( 10'd0 ) : ( n37 ) ;
assign n39 =  ( n16 ) ? ( n38 ) : ( RAM_y ) ;
assign n40 =  ( n25 ) ? ( RAM_y ) : ( RAM_y ) ;
assign n41 =  ( n15 ) ? ( n39 ) : ( n40 ) ;
assign n42 =  ( n12 ) ? ( RAM_y ) : ( n41 ) ;
assign n43 =  ( n6 ) ? ( RAM_y ) : ( n42 ) ;
assign n44 =  ( RAM_x ) > ( 9'd9 )  ;
assign n45 = stencil_8[71:64] ;
assign n46 = stencil_7[71:64] ;
assign n47 = stencil_6[71:64] ;
assign n48 = stencil_5[71:64] ;
assign n49 = stencil_4[71:64] ;
assign n50 = stencil_3[71:64] ;
assign n51 = stencil_2[71:64] ;
assign n52 = stencil_1[71:64] ;
assign n53 = stencil_0[71:64] ;
assign n54 =  { ( n52 ) , ( n53 ) }  ;
assign n55 =  { ( n51 ) , ( n54 ) }  ;
assign n56 =  { ( n50 ) , ( n55 ) }  ;
assign n57 =  { ( n49 ) , ( n56 ) }  ;
assign n58 =  { ( n48 ) , ( n57 ) }  ;
assign n59 =  { ( n47 ) , ( n58 ) }  ;
assign n60 =  { ( n46 ) , ( n59 ) }  ;
assign n61 =  { ( n45 ) , ( n60 ) }  ;
assign n62 = stencil_8[63:56] ;
assign n63 = stencil_7[63:56] ;
assign n64 = stencil_6[63:56] ;
assign n65 = stencil_5[63:56] ;
assign n66 = stencil_4[63:56] ;
assign n67 = stencil_3[63:56] ;
assign n68 = stencil_2[63:56] ;
assign n69 = stencil_1[63:56] ;
assign n70 = stencil_0[63:56] ;
assign n71 =  { ( n69 ) , ( n70 ) }  ;
assign n72 =  { ( n68 ) , ( n71 ) }  ;
assign n73 =  { ( n67 ) , ( n72 ) }  ;
assign n74 =  { ( n66 ) , ( n73 ) }  ;
assign n75 =  { ( n65 ) , ( n74 ) }  ;
assign n76 =  { ( n64 ) , ( n75 ) }  ;
assign n77 =  { ( n63 ) , ( n76 ) }  ;
assign n78 =  { ( n62 ) , ( n77 ) }  ;
assign n79 = stencil_8[55:48] ;
assign n80 = stencil_7[55:48] ;
assign n81 = stencil_6[55:48] ;
assign n82 = stencil_5[55:48] ;
assign n83 = stencil_4[55:48] ;
assign n84 = stencil_3[55:48] ;
assign n85 = stencil_2[55:48] ;
assign n86 = stencil_1[55:48] ;
assign n87 = stencil_0[55:48] ;
assign n88 =  { ( n86 ) , ( n87 ) }  ;
assign n89 =  { ( n85 ) , ( n88 ) }  ;
assign n90 =  { ( n84 ) , ( n89 ) }  ;
assign n91 =  { ( n83 ) , ( n90 ) }  ;
assign n92 =  { ( n82 ) , ( n91 ) }  ;
assign n93 =  { ( n81 ) , ( n92 ) }  ;
assign n94 =  { ( n80 ) , ( n93 ) }  ;
assign n95 =  { ( n79 ) , ( n94 ) }  ;
assign n96 = stencil_8[47:40] ;
assign n97 = stencil_7[47:40] ;
assign n98 = stencil_6[47:40] ;
assign n99 = stencil_5[47:40] ;
assign n100 = stencil_4[47:40] ;
assign n101 = stencil_3[47:40] ;
assign n102 = stencil_2[47:40] ;
assign n103 = stencil_1[47:40] ;
assign n104 = stencil_0[47:40] ;
assign n105 =  { ( n103 ) , ( n104 ) }  ;
assign n106 =  { ( n102 ) , ( n105 ) }  ;
assign n107 =  { ( n101 ) , ( n106 ) }  ;
assign n108 =  { ( n100 ) , ( n107 ) }  ;
assign n109 =  { ( n99 ) , ( n108 ) }  ;
assign n110 =  { ( n98 ) , ( n109 ) }  ;
assign n111 =  { ( n97 ) , ( n110 ) }  ;
assign n112 =  { ( n96 ) , ( n111 ) }  ;
assign n113 = stencil_8[39:32] ;
assign n114 = stencil_7[39:32] ;
assign n115 = stencil_6[39:32] ;
assign n116 = stencil_5[39:32] ;
assign n117 = stencil_4[39:32] ;
assign n118 = stencil_3[39:32] ;
assign n119 = stencil_2[39:32] ;
assign n120 = stencil_1[39:32] ;
assign n121 = stencil_0[39:32] ;
assign n122 =  { ( n120 ) , ( n121 ) }  ;
assign n123 =  { ( n119 ) , ( n122 ) }  ;
assign n124 =  { ( n118 ) , ( n123 ) }  ;
assign n125 =  { ( n117 ) , ( n124 ) }  ;
assign n126 =  { ( n116 ) , ( n125 ) }  ;
assign n127 =  { ( n115 ) , ( n126 ) }  ;
assign n128 =  { ( n114 ) , ( n127 ) }  ;
assign n129 =  { ( n113 ) , ( n128 ) }  ;
assign n130 = stencil_8[31:24] ;
assign n131 = stencil_7[31:24] ;
assign n132 = stencil_6[31:24] ;
assign n133 = stencil_5[31:24] ;
assign n134 = stencil_4[31:24] ;
assign n135 = stencil_3[31:24] ;
assign n136 = stencil_2[31:24] ;
assign n137 = stencil_1[31:24] ;
assign n138 = stencil_0[31:24] ;
assign n139 =  { ( n137 ) , ( n138 ) }  ;
assign n140 =  { ( n136 ) , ( n139 ) }  ;
assign n141 =  { ( n135 ) , ( n140 ) }  ;
assign n142 =  { ( n134 ) , ( n141 ) }  ;
assign n143 =  { ( n133 ) , ( n142 ) }  ;
assign n144 =  { ( n132 ) , ( n143 ) }  ;
assign n145 =  { ( n131 ) , ( n144 ) }  ;
assign n146 =  { ( n130 ) , ( n145 ) }  ;
assign n147 = stencil_8[23:16] ;
assign n148 = stencil_7[23:16] ;
assign n149 = stencil_6[23:16] ;
assign n150 = stencil_5[23:16] ;
assign n151 = stencil_4[23:16] ;
assign n152 = stencil_3[23:16] ;
assign n153 = stencil_2[23:16] ;
assign n154 = stencil_1[23:16] ;
assign n155 = stencil_0[23:16] ;
assign n156 =  { ( n154 ) , ( n155 ) }  ;
assign n157 =  { ( n153 ) , ( n156 ) }  ;
assign n158 =  { ( n152 ) , ( n157 ) }  ;
assign n159 =  { ( n151 ) , ( n158 ) }  ;
assign n160 =  { ( n150 ) , ( n159 ) }  ;
assign n161 =  { ( n149 ) , ( n160 ) }  ;
assign n162 =  { ( n148 ) , ( n161 ) }  ;
assign n163 =  { ( n147 ) , ( n162 ) }  ;
assign n164 = stencil_8[15:8] ;
assign n165 = stencil_7[15:8] ;
assign n166 = stencil_6[15:8] ;
assign n167 = stencil_5[15:8] ;
assign n168 = stencil_4[15:8] ;
assign n169 = stencil_3[15:8] ;
assign n170 = stencil_2[15:8] ;
assign n171 = stencil_1[15:8] ;
assign n172 = stencil_0[15:8] ;
assign n173 =  { ( n171 ) , ( n172 ) }  ;
assign n174 =  { ( n170 ) , ( n173 ) }  ;
assign n175 =  { ( n169 ) , ( n174 ) }  ;
assign n176 =  { ( n168 ) , ( n175 ) }  ;
assign n177 =  { ( n167 ) , ( n176 ) }  ;
assign n178 =  { ( n166 ) , ( n177 ) }  ;
assign n179 =  { ( n165 ) , ( n178 ) }  ;
assign n180 =  { ( n164 ) , ( n179 ) }  ;
assign n181 = stencil_8[7:0] ;
assign n182 = stencil_7[7:0] ;
assign n183 = stencil_6[7:0] ;
assign n184 = stencil_5[7:0] ;
assign n185 = stencil_4[7:0] ;
assign n186 = stencil_3[7:0] ;
assign n187 = stencil_2[7:0] ;
assign n188 = stencil_1[7:0] ;
assign n189 = stencil_0[7:0] ;
assign n190 =  { ( n188 ) , ( n189 ) }  ;
assign n191 =  { ( n187 ) , ( n190 ) }  ;
assign n192 =  { ( n186 ) , ( n191 ) }  ;
assign n193 =  { ( n185 ) , ( n192 ) }  ;
assign n194 =  { ( n184 ) , ( n193 ) }  ;
assign n195 =  { ( n183 ) , ( n194 ) }  ;
assign n196 =  { ( n182 ) , ( n195 ) }  ;
assign n197 =  { ( n181 ) , ( n196 ) }  ;
assign n198 =  { ( n180 ) , ( n197 ) }  ;
assign n199 =  { ( n163 ) , ( n198 ) }  ;
assign n200 =  { ( n146 ) , ( n199 ) }  ;
assign n201 =  { ( n129 ) , ( n200 ) }  ;
assign n202 =  { ( n112 ) , ( n201 ) }  ;
assign n203 =  { ( n95 ) , ( n202 ) }  ;
assign n204 =  { ( n78 ) , ( n203 ) }  ;
assign n205 =  { ( n61 ) , ( n204 ) }  ;
assign n206 =  ( n44 ) ? ( n205 ) : ( proc_in ) ;
assign n207 = gb_fun(n206) ;
assign n208 =  ( n25 ) ? ( arg_0_TDATA ) : ( arg_0_TDATA ) ;
assign n209 =  ( n15 ) ? ( arg_0_TDATA ) : ( n208 ) ;
assign n210 =  ( n12 ) ? ( arg_0_TDATA ) : ( n209 ) ;
assign n211 =  ( n6 ) ? ( n207 ) : ( n210 ) ;
assign n212 =  ( RAM_x ) > ( 9'd8 )  ;
assign n213 =  ( RAM_y ) >= ( 10'd8 )  ;
assign n214 =  ( n212 ) & ( n213 )  ;
assign n215 =  ( RAM_x ) == ( 9'd1 )  ;
assign n216 =  ( RAM_y ) > ( 10'd8 )  ;
assign n217 =  ( n215 ) & ( n216 )  ;
assign n218 =  ( n214 ) | ( n217 )  ;
assign n219 =  ( n218 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n220 =  ( n25 ) ? ( 1'd0 ) : ( arg_0_TVALID ) ;
assign n221 =  ( n15 ) ? ( arg_0_TVALID ) : ( n220 ) ;
assign n222 =  ( n12 ) ? ( 1'd0 ) : ( n221 ) ;
assign n223 =  ( n6 ) ? ( n219 ) : ( n222 ) ;
assign n224 =  ( 10'd648 ) - ( 10'd1 )  ;
assign n225 =  ( RAM_y ) == ( n224 )  ;
assign n226 =  ( n16 ) & ( n225 )  ;
assign n227 =  ( n226 ) ? ( 1'd0 ) : ( 1'd1 ) ;
assign n228 =  ( n226 ) ? ( 1'd1 ) : ( 1'd0 ) ;
assign n229 =  ( n25 ) ? ( 1'd0 ) : ( arg_1_TREADY ) ;
assign n230 =  ( n15 ) ? ( n228 ) : ( n229 ) ;
assign n231 =  ( n12 ) ? ( 1'd1 ) : ( n230 ) ;
assign n232 =  ( n6 ) ? ( n227 ) : ( n231 ) ;
assign n233 =  ( n25 ) ? ( arg_1_TDATA ) : ( cur_pix ) ;
assign n234 =  ( n15 ) ? ( cur_pix ) : ( n233 ) ;
assign n235 =  ( n12 ) ? ( cur_pix ) : ( n234 ) ;
assign n236 =  ( n6 ) ? ( cur_pix ) : ( n235 ) ;
assign n237 =  ( n15 ) ? ( cur_pix ) : ( pre_pix ) ;
assign n238 =  ( n12 ) ? ( cur_pix ) : ( n237 ) ;
assign n239 =  ( n6 ) ? ( pre_pix ) : ( n238 ) ;
assign n240 =  ( n15 ) ? ( proc_in ) : ( proc_in ) ;
assign n241 =  ( n12 ) ? ( proc_in ) : ( n240 ) ;
assign n242 =  ( n6 ) ? ( n206 ) : ( n241 ) ;
assign n243 =  ( n15 ) ? ( n228 ) : ( st_ready ) ;
assign n244 =  ( n12 ) ? ( 1'd1 ) : ( n243 ) ;
assign n245 =  ( n6 ) ? ( 1'd1 ) : ( n244 ) ;
assign n246 =  ( RAM_y ) < ( 10'd8 )  ;
assign n247 =  ( n246 ) ? ( stencil_0 ) : ( stencil_1 ) ;
assign n248 =  ( n25 ) ? ( stencil_0 ) : ( stencil_0 ) ;
assign n249 =  ( n15 ) ? ( stencil_0 ) : ( n248 ) ;
assign n250 =  ( n12 ) ? ( stencil_0 ) : ( n249 ) ;
assign n251 =  ( n6 ) ? ( n247 ) : ( n250 ) ;
assign n252 =  ( n246 ) ? ( stencil_1 ) : ( stencil_2 ) ;
assign n253 =  ( n25 ) ? ( stencil_1 ) : ( stencil_1 ) ;
assign n254 =  ( n15 ) ? ( stencil_1 ) : ( n253 ) ;
assign n255 =  ( n12 ) ? ( stencil_1 ) : ( n254 ) ;
assign n256 =  ( n6 ) ? ( n252 ) : ( n255 ) ;
assign n257 =  ( n246 ) ? ( stencil_2 ) : ( stencil_3 ) ;
assign n258 =  ( n25 ) ? ( stencil_2 ) : ( stencil_2 ) ;
assign n259 =  ( n15 ) ? ( stencil_2 ) : ( n258 ) ;
assign n260 =  ( n12 ) ? ( stencil_2 ) : ( n259 ) ;
assign n261 =  ( n6 ) ? ( n257 ) : ( n260 ) ;
assign n262 =  ( n246 ) ? ( stencil_3 ) : ( stencil_4 ) ;
assign n263 =  ( n25 ) ? ( stencil_3 ) : ( stencil_3 ) ;
assign n264 =  ( n15 ) ? ( stencil_3 ) : ( n263 ) ;
assign n265 =  ( n12 ) ? ( stencil_3 ) : ( n264 ) ;
assign n266 =  ( n6 ) ? ( n262 ) : ( n265 ) ;
assign n267 =  ( n246 ) ? ( stencil_4 ) : ( stencil_5 ) ;
assign n268 =  ( n25 ) ? ( stencil_4 ) : ( stencil_4 ) ;
assign n269 =  ( n15 ) ? ( stencil_4 ) : ( n268 ) ;
assign n270 =  ( n12 ) ? ( stencil_4 ) : ( n269 ) ;
assign n271 =  ( n6 ) ? ( n267 ) : ( n270 ) ;
assign n272 =  ( n246 ) ? ( stencil_5 ) : ( stencil_6 ) ;
assign n273 =  ( n25 ) ? ( stencil_5 ) : ( stencil_5 ) ;
assign n274 =  ( n15 ) ? ( stencil_5 ) : ( n273 ) ;
assign n275 =  ( n12 ) ? ( stencil_5 ) : ( n274 ) ;
assign n276 =  ( n6 ) ? ( n272 ) : ( n275 ) ;
assign n277 =  ( n246 ) ? ( stencil_6 ) : ( stencil_7 ) ;
assign n278 =  ( n25 ) ? ( stencil_6 ) : ( stencil_6 ) ;
assign n279 =  ( n15 ) ? ( stencil_6 ) : ( n278 ) ;
assign n280 =  ( n12 ) ? ( stencil_6 ) : ( n279 ) ;
assign n281 =  ( n6 ) ? ( n277 ) : ( n280 ) ;
assign n282 =  ( n246 ) ? ( stencil_7 ) : ( stencil_8 ) ;
assign n283 =  ( n25 ) ? ( stencil_7 ) : ( stencil_7 ) ;
assign n284 =  ( n15 ) ? ( stencil_7 ) : ( n283 ) ;
assign n285 =  ( n12 ) ? ( stencil_7 ) : ( n284 ) ;
assign n286 =  ( n6 ) ? ( n282 ) : ( n285 ) ;
assign n287 =  ( RAM_w ) == ( 3'd0 )  ;
assign n288 =  ( RAM_x ) - ( 9'd1 )  ;
assign n289 =  (  RAM_7 [ n288 ] )  ;
assign n290 =  ( RAM_w ) == ( 3'd1 )  ;
assign n291 =  ( RAM_w ) == ( 3'd2 )  ;
assign n292 =  ( RAM_w ) == ( 3'd3 )  ;
assign n293 =  ( RAM_w ) == ( 3'd4 )  ;
assign n294 =  ( RAM_w ) == ( 3'd5 )  ;
assign n295 =  ( RAM_w ) == ( 3'd6 )  ;
assign n296 =  (  RAM_6 [ n288 ] )  ;
assign n297 =  ( n295 ) ? ( n289 ) : ( n296 ) ;
assign n298 =  ( n294 ) ? ( n289 ) : ( n297 ) ;
assign n299 =  ( n293 ) ? ( n289 ) : ( n298 ) ;
assign n300 =  ( n292 ) ? ( n289 ) : ( n299 ) ;
assign n301 =  ( n291 ) ? ( n289 ) : ( n300 ) ;
assign n302 =  ( n290 ) ? ( n289 ) : ( n301 ) ;
assign n303 =  ( n287 ) ? ( n289 ) : ( n302 ) ;
assign n304 =  (  RAM_5 [ n288 ] )  ;
assign n305 =  ( n295 ) ? ( n296 ) : ( n304 ) ;
assign n306 =  ( n294 ) ? ( n296 ) : ( n305 ) ;
assign n307 =  ( n293 ) ? ( n296 ) : ( n306 ) ;
assign n308 =  ( n292 ) ? ( n296 ) : ( n307 ) ;
assign n309 =  ( n291 ) ? ( n296 ) : ( n308 ) ;
assign n310 =  ( n290 ) ? ( n296 ) : ( n309 ) ;
assign n311 =  ( n287 ) ? ( n296 ) : ( n310 ) ;
assign n312 =  (  RAM_4 [ n288 ] )  ;
assign n313 =  ( n295 ) ? ( n304 ) : ( n312 ) ;
assign n314 =  ( n294 ) ? ( n304 ) : ( n313 ) ;
assign n315 =  ( n293 ) ? ( n304 ) : ( n314 ) ;
assign n316 =  ( n292 ) ? ( n304 ) : ( n315 ) ;
assign n317 =  ( n291 ) ? ( n304 ) : ( n316 ) ;
assign n318 =  ( n290 ) ? ( n304 ) : ( n317 ) ;
assign n319 =  ( n287 ) ? ( n304 ) : ( n318 ) ;
assign n320 =  (  RAM_3 [ n288 ] )  ;
assign n321 =  ( n295 ) ? ( n312 ) : ( n320 ) ;
assign n322 =  ( n294 ) ? ( n312 ) : ( n321 ) ;
assign n323 =  ( n293 ) ? ( n312 ) : ( n322 ) ;
assign n324 =  ( n292 ) ? ( n312 ) : ( n323 ) ;
assign n325 =  ( n291 ) ? ( n312 ) : ( n324 ) ;
assign n326 =  ( n290 ) ? ( n312 ) : ( n325 ) ;
assign n327 =  ( n287 ) ? ( n312 ) : ( n326 ) ;
assign n328 =  (  RAM_2 [ n288 ] )  ;
assign n329 =  ( n295 ) ? ( n320 ) : ( n328 ) ;
assign n330 =  ( n294 ) ? ( n320 ) : ( n329 ) ;
assign n331 =  ( n293 ) ? ( n320 ) : ( n330 ) ;
assign n332 =  ( n292 ) ? ( n320 ) : ( n331 ) ;
assign n333 =  ( n291 ) ? ( n320 ) : ( n332 ) ;
assign n334 =  ( n290 ) ? ( n320 ) : ( n333 ) ;
assign n335 =  ( n287 ) ? ( n320 ) : ( n334 ) ;
assign n336 =  (  RAM_1 [ n288 ] )  ;
assign n337 =  ( n295 ) ? ( n328 ) : ( n336 ) ;
assign n338 =  ( n294 ) ? ( n328 ) : ( n337 ) ;
assign n339 =  ( n293 ) ? ( n328 ) : ( n338 ) ;
assign n340 =  ( n292 ) ? ( n328 ) : ( n339 ) ;
assign n341 =  ( n291 ) ? ( n328 ) : ( n340 ) ;
assign n342 =  ( n290 ) ? ( n328 ) : ( n341 ) ;
assign n343 =  ( n287 ) ? ( n328 ) : ( n342 ) ;
assign n344 =  (  RAM_0 [ n288 ] )  ;
assign n345 =  ( n295 ) ? ( n336 ) : ( n344 ) ;
assign n346 =  ( n294 ) ? ( n336 ) : ( n345 ) ;
assign n347 =  ( n293 ) ? ( n336 ) : ( n346 ) ;
assign n348 =  ( n292 ) ? ( n336 ) : ( n347 ) ;
assign n349 =  ( n291 ) ? ( n336 ) : ( n348 ) ;
assign n350 =  ( n290 ) ? ( n336 ) : ( n349 ) ;
assign n351 =  ( n287 ) ? ( n336 ) : ( n350 ) ;
assign n352 =  ( n295 ) ? ( n344 ) : ( n289 ) ;
assign n353 =  ( n294 ) ? ( n344 ) : ( n352 ) ;
assign n354 =  ( n293 ) ? ( n344 ) : ( n353 ) ;
assign n355 =  ( n292 ) ? ( n344 ) : ( n354 ) ;
assign n356 =  ( n291 ) ? ( n344 ) : ( n355 ) ;
assign n357 =  ( n290 ) ? ( n344 ) : ( n356 ) ;
assign n358 =  ( n287 ) ? ( n344 ) : ( n357 ) ;
assign n359 =  { ( n351 ) , ( n358 ) }  ;
assign n360 =  { ( n343 ) , ( n359 ) }  ;
assign n361 =  { ( n335 ) , ( n360 ) }  ;
assign n362 =  { ( n327 ) , ( n361 ) }  ;
assign n363 =  { ( n319 ) , ( n362 ) }  ;
assign n364 =  { ( n311 ) , ( n363 ) }  ;
assign n365 =  { ( n303 ) , ( n364 ) }  ;
assign n366 =  { ( pre_pix ) , ( n365 ) }  ;
assign n367 =  ( n246 ) ? ( stencil_8 ) : ( n366 ) ;
assign n368 =  ( n25 ) ? ( stencil_8 ) : ( stencil_8 ) ;
assign n369 =  ( n15 ) ? ( n367 ) : ( n368 ) ;
assign n370 =  ( n12 ) ? ( stencil_8 ) : ( n369 ) ;
assign n371 =  ( n6 ) ? ( stencil_8 ) : ( n370 ) ;
assign n372 = ~ ( n6 ) ;
assign n373 = ~ ( n12 ) ;
assign n374 =  ( n372 ) & ( n373 )  ;
assign n375 = ~ ( n15 ) ;
assign n376 =  ( n374 ) & ( n375 )  ;
assign n377 = ~ ( n25 ) ;
assign n378 =  ( n376 ) & ( n377 )  ;
assign n379 =  ( n376 ) & ( n25 )  ;
assign n380 =  ( n374 ) & ( n15 )  ;
assign n381 = ~ ( n287 ) ;
assign n382 =  ( n380 ) & ( n381 )  ;
assign n383 =  ( n380 ) & ( n287 )  ;
assign n384 =  ( n372 ) & ( n12 )  ;
assign RAM_0_addr0 = n383 ? (n288) : (0);
assign RAM_0_data0 = n383 ? (pre_pix) : (RAM_0[0]);
assign n385 = ~ ( n290 ) ;
assign n386 =  ( n380 ) & ( n385 )  ;
assign n387 =  ( n380 ) & ( n290 )  ;
assign RAM_1_addr0 = n387 ? (n288) : (0);
assign RAM_1_data0 = n387 ? (pre_pix) : (RAM_1[0]);
assign n388 = ~ ( n291 ) ;
assign n389 =  ( n380 ) & ( n388 )  ;
assign n390 =  ( n380 ) & ( n291 )  ;
assign RAM_2_addr0 = n390 ? (n288) : (0);
assign RAM_2_data0 = n390 ? (pre_pix) : (RAM_2[0]);
assign n391 = ~ ( n292 ) ;
assign n392 =  ( n380 ) & ( n391 )  ;
assign n393 =  ( n380 ) & ( n292 )  ;
assign RAM_3_addr0 = n393 ? (n288) : (0);
assign RAM_3_data0 = n393 ? (pre_pix) : (RAM_3[0]);
assign n394 = ~ ( n293 ) ;
assign n395 =  ( n380 ) & ( n394 )  ;
assign n396 =  ( n380 ) & ( n293 )  ;
assign RAM_4_addr0 = n396 ? (n288) : (0);
assign RAM_4_data0 = n396 ? (pre_pix) : (RAM_4[0]);
assign n397 = ~ ( n294 ) ;
assign n398 =  ( n380 ) & ( n397 )  ;
assign n399 =  ( n380 ) & ( n294 )  ;
assign RAM_5_addr0 = n399 ? (n288) : (0);
assign RAM_5_data0 = n399 ? (pre_pix) : (RAM_5[0]);
assign n400 = ~ ( n295 ) ;
assign n401 =  ( n380 ) & ( n400 )  ;
assign n402 =  ( n380 ) & ( n295 )  ;
assign RAM_6_addr0 = n402 ? (n288) : (0);
assign RAM_6_data0 = n402 ? (pre_pix) : (RAM_6[0]);
assign n403 = ~ ( n17 ) ;
assign n404 =  ( n380 ) & ( n403 )  ;
assign n405 =  ( n380 ) & ( n17 )  ;
assign RAM_7_addr0 = n405 ? (n288) : (0);
assign RAM_7_data0 = n405 ? (pre_pix) : (RAM_7[0]);
function [7:0] gb_fun ;
input [647:0] arg0;
    begin
//TODO: Add the specific function HERE.    end
endfunction

always @(posedge clk) begin
   if(rst) begin
       RAM_w <= RAM_w;
       RAM_x <= RAM_x;
       RAM_y <= RAM_y;
       arg_0_TDATA <= arg_0_TDATA;
       arg_0_TVALID <= arg_0_TVALID;
       arg_1_TREADY <= arg_1_TREADY;
       cur_pix <= cur_pix;
       pre_pix <= pre_pix;
       proc_in <= proc_in;
       st_ready <= st_ready;
       stencil_0 <= stencil_0;
       stencil_1 <= stencil_1;
       stencil_2 <= stencil_2;
       stencil_3 <= stencil_3;
       stencil_4 <= stencil_4;
       stencil_5 <= stencil_5;
       stencil_6 <= stencil_6;
       stencil_7 <= stencil_7;
       stencil_8 <= stencil_8;
   end
   else if(step) begin
       RAM_w <= n29;
       RAM_x <= n35;
       RAM_y <= n43;
       arg_0_TDATA <= n211;
       arg_0_TVALID <= n223;
       arg_1_TREADY <= n232;
       cur_pix <= n236;
       pre_pix <= n239;
       proc_in <= n242;
       st_ready <= n245;
       stencil_0 <= n251;
       stencil_1 <= n256;
       stencil_2 <= n261;
       stencil_3 <= n266;
       stencil_4 <= n271;
       stencil_5 <= n276;
       stencil_6 <= n281;
       stencil_7 <= n286;
       stencil_8 <= n371;
       RAM_0 [ RAM_0_addr0 ] <= RAM_0_data0;
       RAM_1 [ RAM_1_addr0 ] <= RAM_1_data0;
       RAM_2 [ RAM_2_addr0 ] <= RAM_2_data0;
       RAM_3 [ RAM_3_addr0 ] <= RAM_3_data0;
       RAM_4 [ RAM_4_addr0 ] <= RAM_4_data0;
       RAM_5 [ RAM_5_addr0 ] <= RAM_5_data0;
       RAM_6 [ RAM_6_addr0 ] <= RAM_6_data0;
       RAM_7 [ RAM_7_addr0 ] <= RAM_7_data0;
   end
end
endmodule
